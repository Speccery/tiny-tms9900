//
// Simplistic 4096x16 RAM module
//
// This source code is public domain
//

module ROM(CLK, nCS, ADDR, DO);

  // Port definition
  input CLK, nCS;
  input  [11:0] ADDR;
  output [15:0] DO;
  
  wire          CLK, nCS;
  wire   [11:0] ADDR;
  reg    [15:0] DO;
  
  // Implementation
  reg [15:0] mem[4095:0];
  
  always @(posedge CLK)
  begin
    if (!nCS) begin
      DO = mem[ADDR];
    end
  end
  
  initial
  begin
    mem[0000]='hec00; mem[0001]='h0226; mem[0002]='hf0d6; mem[0003]='hf0f6; mem[0004]='hf0ca; mem[0005]='hf0ea; mem[0006]='hf0be; mem[0007]='hf0de; // address 0x0000
    mem[0008]='hf0b2; mem[0009]='hf0d2; mem[0010]='h0d0a; mem[0011]='h4d4f; mem[0012]='h4e3f; mem[0013]='h2000; mem[0014]='h2020; mem[0015]='h2020; // address 0x0010
    mem[0016]='h2020; mem[0017]='h000d; mem[0018]='h0a42; mem[0019]='h5000; mem[0020]='h4944; mem[0021]='h543d; mem[0022]='h000d; mem[0023]='h0a52; // address 0x0020
    mem[0024]='h4541; mem[0025]='h4459; mem[0026]='h2059; mem[0027]='h2f4e; mem[0028]='h2000; mem[0029]='h5700; mem[0030]='h5000; mem[0031]='h5300; // address 0x0030
    mem[0032]='hf0ac; mem[0033]='hf0be; mem[0034]='hf09e; mem[0035]='hf0b0; mem[0036]='hf090; mem[0037]='hf0a2; mem[0038]='hf082; mem[0039]='hf094; // address 0x0040
    mem[0040]='hf074; mem[0041]='hf086; mem[0042]='hf066; mem[0043]='hf078; mem[0044]='hf058; mem[0045]='hf06a; mem[0046]='hf04a; mem[0047]='hf05c; // address 0x0050
    mem[0048]='hec24; mem[0049]='h03f8; mem[0050]='hec24; mem[0051]='h0396; mem[0052]='hec24; mem[0053]='h0402; mem[0054]='hec0a; mem[0055]='h0326; // address 0x0060
    mem[0056]='hec16; mem[0057]='h02ee; mem[0058]='hec16; mem[0059]='h02e2; mem[0060]='hec24; mem[0061]='h032c; mem[0062]='hec00; mem[0063]='h0442; // address 0x0070

// trying with these settings:
    mem[0064]='h0460; mem[0065]='h0142; 
    
    // Bitrate table in the original ROM
    mem[0066]='h0009; mem[0067]='h0034;   // First word is some count, second the value to write to TMS9902
    mem[0068]='h0012; mem[0069]='h0034; 
    mem[0070]='h0023; mem[0071]='h0034; // address 0x0080
    mem[0072]='h0046; mem[0073]='h0034; 
    mem[0074]='h008d; mem[0075]='h0034; 
    mem[0076]='h0119; mem[0077]='h0034; 
    mem[0078]='h02a4; mem[0079]='h0034; // address 0x0090
    mem[0080]='h7fff; mem[0081]='h0034; 
    
    mem[0082]='h0d0a; mem[0083]='h4552; mem[0084]='h524f; mem[0085]='h5220; mem[0086]='h000d; mem[0087]='h0a45; // address 0x00a0


// In the verilog simulation environment I had these lines
//    mem[0064]='h0460; mem[0065]='h0142; mem[0066]='h0009; mem[0067]='h0001; mem[0068]='h0012; mem[0069]='h0001; mem[0070]='h0023; mem[0071]='h0001; // address 0x0080
//    mem[0072]='h0046; mem[0073]='h0001; mem[0074]='h008d; mem[0075]='h0001; mem[0076]='h0119; mem[0077]='h0001; mem[0078]='h02a4; mem[0079]='h0001; // address 0x0090
//    mem[0080]='h7fff; mem[0081]='h0001; mem[0082]='h0d0a; mem[0083]='h4552; mem[0084]='h524f; mem[0085]='h5220; mem[0086]='h000d; mem[0087]='h0a45; // address 0x00a0
  
// this used to be commented out
//  mem[0064]='h0460; mem[0065]='h0142; mem[0066]='h0009; mem[0067]='h001a; mem[0068]='h0012; mem[0069]='h0034; mem[0070]='h0023; mem[0071]='h0068; // address 0x0080
//  mem[0072]='h0046; mem[0073]='h00d0; mem[0074]='h008d; mem[0075]='h01a1; mem[0076]='h0119; mem[0077]='h0341; mem[0078]='h02a4; mem[0079]='h04d0; // address 0x0090
//  mem[0080]='h7fff; mem[0081]='h0638; mem[0082]='h0d0a; mem[0083]='h4552; mem[0084]='h524f; mem[0085]='h5220; mem[0086]='h000d; mem[0087]='h0a45; // address 0x00a0

    mem[0088]='h564d; mem[0089]='h4255; mem[0090]='h4720; mem[0091]='h2052; mem[0092]='h312e; mem[0093]='h3000; mem[0094]='h0d0a; mem[0095]='h5200; // address 0x00b0
    mem[0096]='h0d0a; mem[0097]='h4831; mem[0098]='h2b48; mem[0099]='h323d; mem[0100]='h0020; mem[0101]='h4831; mem[0102]='h2d48; mem[0103]='h323d; // address 0x00c0
    mem[0104]='h0020; mem[0105]='h4552; mem[0106]='h524f; mem[0107]='h5200; mem[0108]='h0d0a; mem[0109]='h434f; mem[0110]='h4d3f; mem[0111]='h2000; // address 0x00d0
    mem[0112]='h3a0d; mem[0113]='h000d; mem[0114]='h0a54; mem[0115]='h4552; mem[0116]='h4d49; mem[0117]='h4e41; mem[0118]='h4c20; mem[0119]='h4d4f; // address 0x00e0
    mem[0120]='h4445; mem[0121]='h0d0a; mem[0122]='h000d; mem[0123]='h0a43; mem[0124]='h4d44; mem[0125]='h2045; mem[0126]='h5252; mem[0127]='h000d; // address 0x00f0
    mem[0128]='h0a50; mem[0129]='h4152; mem[0130]='h4d20; mem[0131]='h4552; mem[0132]='h5200; mem[0133]='h0d0a; mem[0134]='h434b; mem[0135]='h534d; // address 0x0100
    mem[0136]='h2045; mem[0137]='h5252; mem[0138]='h000d; mem[0139]='h0a54; mem[0140]='h4147; mem[0141]='h2045; mem[0142]='h5252; mem[0143]='h0055; // address 0x0110
    mem[0144]='h504c; mem[0145]='h4420; mem[0146]='h4552; mem[0147]='h5200; mem[0148]='h460d; mem[0149]='h000a; mem[0150]='h7f3a; mem[0151]='h0d0a; // address 0x0120
    mem[0152]='h7f13; mem[0153]='h0d14; mem[0154]='h7f00; mem[0155]='h120a; mem[0156]='h7f00; 
    
    // Here at 157 (013A) we have the configuration bytes; the default word is 'h6242
    // mem[0157]='h6242; 
    // 62 = (0110 0010) 7 bits/character, even parity, 2 stop bits.
    // 42 = (0100 0010) 7 bits/character, no parity, 2 stop bits.
    // My calculation is that 83 (hex) wound be 8N1
    mem[0157]='h8383; 
    
    mem[0158]='h1100; mem[0159]='h0000; // address 0x0130
    mem[0160]='h0400; mem[0161]='h02e0; mem[0162]='hec00; mem[0163]='h04c1; mem[0164]='h0202; mem[0165]='hfffc; mem[0166]='hccb1; mem[0167]='h0201; // address 0x0140
    mem[0168]='h042e; mem[0169]='hcc81; mem[0170]='h0209; mem[0171]='h0142; mem[0172]='h04c1; mem[0173]='h0641; mem[0174]='h13fe; mem[0175]='hc320; // address 0x0150
    mem[0176]='h013e; mem[0177]='hc80c; mem[0178]='hec2e; mem[0179]='h1f15; mem[0180]='h1601; mem[0181]='h2f45; mem[0182]='h2fa0; mem[0183]='h0014; // address 0x0160
    mem[0184]='h04c0; mem[0185]='h0202; mem[0186]='h0a05; mem[0187]='h0203; mem[0188]='h0004; mem[0189]='h04c4; mem[0190]='h0208; mem[0191]='h0001; // address 0x0170
    mem[0192]='h2ec5; mem[0193]='h0285; mem[0194]='h0d00; mem[0195]='h1604; mem[0196]='h0205; mem[0197]='h0a00; mem[0198]='h2f05; mem[0199]='h1019; // address 0x0180
    mem[0200]='h0285; mem[0201]='h2000; mem[0202]='h1316; mem[0203]='h0285; mem[0204]='h2c00; mem[0205]='h1313; mem[0206]='h0285; mem[0207]='h4100; // address 0x0190
    mem[0208]='h113c; mem[0209]='h0285; mem[0210]='h5a00; mem[0211]='h1539; mem[0212]='h0603; mem[0213]='h1337; mem[0214]='h06c5; mem[0215]='h0245; // address 0x01a0
    mem[0216]='h001f; mem[0217]='h0283; mem[0218]='h0003; mem[0219]='h1301; mem[0220]='h0482; mem[0221]='ha105; mem[0222]='h0222; mem[0223]='h0050; // address 0x01b0
    mem[0224]='h10df; mem[0225]='h020b; mem[0226]='h027a; mem[0227]='h1002; mem[0228]='h022b; mem[0229]='h0004; mem[0230]='hc2bb; mem[0231]='h1325; // address 0x01c0
    mem[0232]='h810a; mem[0233]='h16fa; mem[0234]='hc1bb; mem[0235]='hc2db; mem[0236]='h0207; mem[0237]='hec00; mem[0238]='h0285; mem[0239]='h0a00; // address 0x01d0
    mem[0240]='h130f; mem[0241]='h0916; mem[0242]='h170e; mem[0243]='h2e44; mem[0244]='h01f8; mem[0245]='h020e; mem[0246]='hcdc4; mem[0247]='h0583; // address 0x01e0
    mem[0248]='h0285; mem[0249]='h0d00; mem[0250]='h1306; mem[0251]='h10f5; mem[0252]='h05c7; mem[0253]='h0285; mem[0254]='h0d00; mem[0255]='h16f7; // address 0x01f0
    mem[0256]='h04c3; mem[0257]='h045b; mem[0258]='h04c0; mem[0259]='h100b; mem[0260]='h0200; mem[0261]='h0001; mem[0262]='h1008; mem[0263]='h0200; // address 0x0200
    mem[0264]='h0002; mem[0265]='h1005; mem[0266]='h0200; mem[0267]='h0003; mem[0268]='h1002; mem[0269]='h0200; mem[0270]='h0004; mem[0271]='h2fa0; // address 0x0210
    mem[0272]='h00a4; mem[0273]='h2e00; mem[0274]='h108e; mem[0275]='h020c; mem[0276]='hec44; mem[0277]='h04fc; mem[0278]='h073c; mem[0279]='h04fc; // address 0x0220
    mem[0280]='h04dc; mem[0281]='hc320; mem[0282]='h013e; mem[0283]='hc80c; mem[0284]='hec2e; mem[0285]='h1d1f; mem[0286]='h04c3; mem[0287]='h3220; // address 0x0230
    mem[0288]='h013a; mem[0289]='h1e0d; mem[0290]='h1f0f; mem[0291]='h13fe; mem[0292]='h0583; mem[0293]='h1f0f; mem[0294]='h16fd; mem[0295]='h0207; // address 0x0240
    mem[0296]='h0084; mem[0297]='h8dc3; mem[0298]='h1102; mem[0299]='h05c7; mem[0300]='h10fc; mem[0301]='h3317; mem[0302]='hc1d7; mem[0303]='h0287; // address 0x0250
    mem[0304]='h01a1; mem[0305]='h1108; mem[0306]='h1602; mem[0307]='h0720; mem[0308]='hec44; mem[0309]='h2f45; mem[0310]='h2fa0; mem[0311]='h00ad; // address 0x0260
    mem[0312]='h0460; mem[0313]='h0142; mem[0314]='h05a0; mem[0315]='hec44; mem[0316]='h10f8; mem[0317]='h01a9; mem[0318]='h0001; mem[0319]='h036c; // address 0x0270
    mem[0320]='h01a4; mem[0321]='h0003; mem[0322]='h0334; mem[0323]='h4ae9; mem[0324]='h0001; mem[0325]='h04ac; mem[0326]='h0305; mem[0327]='h0000; // address 0x0280
    mem[0328]='h042c; mem[0329]='h0b05; mem[0330]='h0001; mem[0331]='h0436; mem[0332]='h0273; mem[0333]='h0000; mem[0334]='h0426; mem[0335]='h0dac; // address 0x0290
    mem[0336]='h0001; mem[0337]='h064a; mem[0338]='h0da4; mem[0339]='h0007; mem[0340]='h0552; mem[0341]='h0069; mem[0342]='h0003; mem[0343]='h0460; // address 0x02a0
    mem[0344]='h0249; mem[0345]='h0000; mem[0346]='h051a; mem[0347]='h0086; mem[0348]='h0007; mem[0349]='h0770; mem[0350]='h60a8; mem[0351]='h0003; // address 0x02b0
    mem[0352]='h07a0; mem[0353]='h19d4; mem[0354]='h0000; mem[0355]='h07b4; mem[0356]='h1438; mem[0357]='h0001; mem[0358]='h07c2; mem[0359]='h0038; // address 0x02c0
    mem[0360]='h0001; mem[0361]='h07ba; mem[0362]='h3078; mem[0363]='h0000; mem[0364]='h0e1a; mem[0365]='h0658; mem[0366]='h0003; mem[0367]='h1166; // address 0x02d0
    mem[0368]='h0000; mem[0369]='h1f15; mem[0370]='h16fe; mem[0371]='h04db; mem[0372]='h361b; mem[0373]='h1e12; mem[0374]='h0380; mem[0375]='h020a; // address 0x02e0
    mem[0376]='h186a; mem[0377]='h1d10; mem[0378]='h1f16; mem[0379]='h16fe; mem[0380]='h321b; mem[0381]='hd2db; mem[0382]='h980b; mem[0383]='h00f2; // address 0x02f0
    mem[0384]='h160b; mem[0385]='hc2e0; mem[0386]='hec44; mem[0387]='h150e; mem[0388]='h0a3a; mem[0389]='h1f16; mem[0390]='h16fe; mem[0391]='h1f17; // address 0x0300
    mem[0392]='h16fc; mem[0393]='h060a; mem[0394]='h16fe; mem[0395]='h0380; mem[0396]='hc2e0; mem[0397]='hec46; mem[0398]='h1303; mem[0399]='hc2e0; // address 0x0310
    mem[0400]='hec44; mem[0401]='h11f3; mem[0402]='h0380; mem[0403]='h2f5b; mem[0404]='h2f1b; mem[0405]='h0380; mem[0406]='hd33b; mem[0407]='h13fd; // address 0x0320
    mem[0408]='h2f0c; mem[0409]='h10fc; mem[0410]='h4008; mem[0411]='h4048; mem[0412]='h0203; mem[0413]='h0008; mem[0414]='h2fa0; mem[0415]='h00f2; // address 0x0330
    mem[0416]='h2e80; mem[0417]='h2fa0; mem[0418]='h00cf; mem[0419]='h2e90; mem[0420]='h1f15; mem[0421]='h1602; mem[0422]='h2f40; mem[0423]='h0459; // address 0x0340
    mem[0424]='h8040; mem[0425]='h13fd; mem[0426]='h05c0; mem[0427]='h0603; mem[0428]='h0283; mem[0429]='h0004; mem[0430]='h1602; mem[0431]='h2fa0; // address 0x0350
    mem[0432]='h0020; mem[0433]='hc0c3; mem[0434]='h13e9; mem[0435]='h2fa0; mem[0436]='h0020; mem[0437]='h10ed; mem[0438]='h4008; mem[0439]='h1004; // address 0x0360
    mem[0440]='h0640; mem[0441]='h0a25; mem[0442]='h16fb; mem[0443]='h8c30; mem[0444]='h2fa0; mem[0445]='h00f2; mem[0446]='h2e80; mem[0447]='h2fa0; // address 0x0370
    mem[0448]='h00cf; mem[0449]='h2e90; mem[0450]='h2fa0; mem[0451]='h0020; mem[0452]='h2e44; mem[0453]='h0390; mem[0454]='h020e; mem[0455]='hc404; // address 0x0380
    mem[0456]='h0a25; mem[0457]='h11ee; mem[0458]='h0459; mem[0459]='h04c9; mem[0460]='h04cc; mem[0461]='h2eca; mem[0462]='h028a; mem[0463]='h3000; // address 0x0390
    mem[0464]='h1a11; mem[0465]='h028a; mem[0466]='h3900; mem[0467]='h1208; mem[0468]='h028a; mem[0469]='h4100; mem[0470]='h1a0b; mem[0471]='h028a; // address 0x03a0
    mem[0472]='h4600; mem[0473]='h1b08; mem[0474]='h022a; mem[0475]='h0900; mem[0476]='h0a4a; mem[0477]='h09ca; mem[0478]='h0a4c; mem[0479]='ha30a; // address 0x03b0
    mem[0480]='h0589; mem[0481]='h10eb; mem[0482]='h028a; mem[0483]='h2000; mem[0484]='h130b; mem[0485]='h028a; mem[0486]='h2d00; mem[0487]='h1308; // address 0x03c0
    mem[0488]='h028a; mem[0489]='h0d00; mem[0490]='h1305; mem[0491]='h028a; mem[0492]='h2c00; mem[0493]='h160c; mem[0494]='h020a; mem[0495]='h2000; // address 0x03d0
    mem[0496]='hc249; mem[0497]='h1304; mem[0498]='hcecc; mem[0499]='hc6ca; mem[0500]='h8fbe; mem[0501]='h0380; mem[0502]='h05cb; mem[0503]='hc6ca; // address 0x03e0
    mem[0504]='hc39e; mem[0505]='h0380; mem[0506]='h05ce; mem[0507]='h10fc; mem[0508]='hc31b; mem[0509]='h0acc; mem[0510]='h0209; mem[0511]='h0001; // address 0x03f0
    mem[0512]='h1003; mem[0513]='hc31b; mem[0514]='h0209; mem[0515]='h0004; mem[0516]='hc28c; mem[0517]='h09ca; mem[0518]='h0a8a; mem[0519]='h028a; // address 0x0400
    mem[0520]='h0900; mem[0521]='h1202; mem[0522]='h022a; mem[0523]='h0700; mem[0524]='h022a; mem[0525]='h3000; mem[0526]='h2f0a; mem[0527]='h0bcc; // address 0x0410
    mem[0528]='h0609; mem[0529]='h16f2; mem[0530]='h0380; mem[0531]='h0207; mem[0532]='h9900; mem[0533]='h03e0; mem[0534]='h0380; mem[0535]='h0287; // address 0x0420
    mem[0536]='h9900; mem[0537]='h130b; mem[0538]='h1013; mem[0539]='h4008; mem[0540]='hc190; mem[0541]='hc420; mem[0542]='h0440; mem[0543]='h0380; // address 0x0430
    mem[0544]='h2fc0; mem[0545]='h064e; mem[0546]='hc406; mem[0547]='h2fa0; mem[0548]='h0023; mem[0549]='h04c7; mem[0550]='h020a; mem[0551]='hfffa; // address 0x0440
    mem[0552]='h2fa0; mem[0553]='h001e; mem[0554]='h2eaa; mem[0555]='hec20; mem[0556]='h05ca; mem[0557]='h16fa; mem[0558]='h0460; mem[0559]='h0142; // address 0x0450
    mem[0560]='hc300; mem[0561]='h04c7; mem[0562]='h0241; mem[0563]='h000f; mem[0564]='h1303; mem[0565]='h0281; mem[0566]='h0009; mem[0567]='h1a01; // address 0x0460
    mem[0568]='h0587; mem[0569]='h0a61; mem[0570]='h0208; mem[0571]='h3406; mem[0572]='he201; mem[0573]='h0488; mem[0574]='h2fa0; mem[0575]='h00f2; // address 0x0470
    mem[0576]='h2e8c; mem[0577]='h2fa0; mem[0578]='h00cf; mem[0579]='hc1c7; mem[0580]='h1601; mem[0581]='h0986; mem[0582]='h2e86; mem[0583]='h2fa0; // address 0x0480
    mem[0584]='h0020; mem[0585]='h2e44; mem[0586]='h04a6; mem[0587]='h020e; mem[0588]='hc184; mem[0589]='hc1c7; mem[0590]='h1601; mem[0591]='h0a86; // address 0x0490
    mem[0592]='h0248; mem[0593]='hf3ff; mem[0594]='h0488; mem[0595]='h09c5; mem[0596]='h16e5; mem[0597]='h0459; mem[0598]='hc1cd; mem[0599]='hc0c3; // address 0x04a0
    mem[0600]='h131f; mem[0601]='h0240; mem[0602]='h000f; mem[0603]='hc180; mem[0604]='h0a10; mem[0605]='ha1c0; mem[0606]='h2fa0; mem[0607]='h00bc; // address 0x04b0
    mem[0608]='h2e06; mem[0609]='h2fa0; mem[0610]='h00cf; mem[0611]='h2e97; mem[0612]='h2fa0; mem[0613]='h0020; mem[0614]='h2e44; mem[0615]='h04d4; // address 0x04c0
    mem[0616]='h020e; mem[0617]='hc5c4; mem[0618]='h0a25; mem[0619]='h153c; mem[0620]='h0a15; mem[0621]='h1304; mem[0622]='h0606; mem[0623]='h1138; // address 0x04d0
    mem[0624]='h0647; mem[0625]='h10ec; mem[0626]='h0286; mem[0627]='h000f; mem[0628]='h1333; mem[0629]='h0586; mem[0630]='h05c7; mem[0631]='h10e6; // address 0x04e0
    mem[0632]='h04c6; mem[0633]='hc1cd; mem[0634]='h2fa0; mem[0635]='h00bc; mem[0636]='h2e06; mem[0637]='h2fa0; mem[0638]='h00cf; mem[0639]='h2e97; // address 0x04f0
    mem[0640]='h0586; mem[0641]='h05c7; mem[0642]='h0286; mem[0643]='h0008; mem[0644]='h13f5; mem[0645]='h0286; mem[0646]='h0010; mem[0647]='h1320; // address 0x0500
    mem[0648]='h2fa0; mem[0649]='h0020; mem[0650]='h2fa0; mem[0651]='h00d6; mem[0652]='h10ef; mem[0653]='h0206; mem[0654]='h003a; mem[0655]='h0207; // address 0x0510
    mem[0656]='h0003; mem[0657]='h0208; mem[0658]='hec1a; mem[0659]='h2fa0; mem[0660]='h00f2; mem[0661]='h2f96; mem[0662]='h2fa0; mem[0663]='h00cf; // address 0x0520
    mem[0664]='hc118; mem[0665]='h2e98; mem[0666]='h2fa0; mem[0667]='h0020; mem[0668]='h2e44; mem[0669]='h053e; mem[0670]='h020e; mem[0671]='hc604; // address 0x0530
    mem[0672]='h0a25; mem[0673]='h1506; mem[0674]='h0a15; mem[0675]='h16ef; mem[0676]='h05c6; mem[0677]='h05c8; mem[0678]='h0607; mem[0679]='h16eb; // address 0x0540
    mem[0680]='h0459; mem[0681]='h4008; mem[0682]='h4048; mem[0683]='h4088; mem[0684]='h8040; mem[0685]='h1202; mem[0686]='h0460; mem[0687]='h0214; // address 0x0550
    mem[0688]='h04c4; mem[0689]='h04c3; mem[0690]='h2fa0; mem[0691]='h0028; mem[0692]='h2f44; mem[0693]='h0284; mem[0694]='h0d00; mem[0695]='h1603; // address 0x0560
    mem[0696]='h0204; mem[0697]='h2000; mem[0698]='h1001; mem[0699]='h2f04; mem[0700]='hd8c4; mem[0701]='hec0c; mem[0702]='h0583; mem[0703]='h0283; // address 0x0570
    mem[0704]='h0008; mem[0705]='h1304; mem[0706]='h0284; mem[0707]='h2000; mem[0708]='h16ef; mem[0709]='h10f6; mem[0710]='h2fa0; mem[0711]='h002d; // address 0x0580
    mem[0712]='h2f44; mem[0713]='h0284; mem[0714]='h5900; mem[0715]='h1641; mem[0716]='h04e0; mem[0717]='hec46; mem[0718]='h2fa0; mem[0719]='h0136; // address 0x0590
    mem[0720]='h04ca; mem[0721]='h04c5; mem[0722]='h06a0; mem[0723]='h061c; mem[0724]='h3000; mem[0725]='h2fa0; mem[0726]='hec0c; mem[0727]='h0203; // address 0x05a0
    mem[0728]='h0008; mem[0729]='hd123; mem[0730]='hec0b; mem[0731]='h0984; mem[0732]='ha144; mem[0733]='h0603; mem[0734]='h16fa; mem[0735]='hc282; // address 0x05b0
    mem[0736]='h06a0; mem[0737]='h061c; mem[0738]='h3100; mem[0739]='hc280; mem[0740]='h06a0; mem[0741]='h061c; mem[0742]='h3900; mem[0743]='hc290; // address 0x05c0
    mem[0744]='h06a0; mem[0745]='h061c; mem[0746]='h4200; mem[0747]='h8040; mem[0748]='h1304; mem[0749]='h05c0; mem[0750]='h0283; mem[0751]='h003c; // address 0x05d0
    mem[0752]='h1af6; mem[0753]='h0225; mem[0754]='h0037; mem[0755]='hc285; mem[0756]='h050a; mem[0757]='h06a0; mem[0758]='h061c; mem[0759]='h3700; // address 0x05e0
    mem[0760]='h04c5; mem[0761]='h2fa0; mem[0762]='h0128; mem[0763]='h8040; mem[0764]='h1304; mem[0765]='h04c3; mem[0766]='h2fa0; mem[0767]='h0137; // address 0x05f0
    mem[0768]='h10e2; mem[0769]='h2fa0; mem[0770]='h012b; mem[0771]='h0203; mem[0772]='h003c; mem[0773]='h2fa0; mem[0774]='h0134; mem[0775]='h0603; // address 0x0600
    mem[0776]='h16fc; mem[0777]='h0720; mem[0778]='hec46; mem[0779]='h2fa0; mem[0780]='h00f2; mem[0781]='h104a; mem[0782]='hc13b; mem[0783]='h2f04; // address 0x0610
    mem[0784]='h0984; mem[0785]='ha144; mem[0786]='h2e8a; mem[0787]='h0223; mem[0788]='h0005; mem[0789]='h0204; mem[0790]='h0004; mem[0791]='h0b4a; // address 0x0620
    mem[0792]='hc30a; mem[0793]='h09cc; mem[0794]='ha14c; mem[0795]='h0225; mem[0796]='h0030; mem[0797]='h028c; mem[0798]='h000a; mem[0799]='h1a02; // address 0x0630
    mem[0800]='h0225; mem[0801]='h0007; mem[0802]='h0604; mem[0803]='h16f3; mem[0804]='h045b; mem[0805]='h2fa0; mem[0806]='h002d; mem[0807]='h2f44; // address 0x0640
    mem[0808]='h0284; mem[0809]='h5900; mem[0810]='h162d; mem[0811]='h0206; mem[0812]='h1100; mem[0813]='h2f06; mem[0814]='h04c7; mem[0815]='h04c8; // address 0x0650
    mem[0816]='h06a0; mem[0817]='h0728; mem[0818]='h100b; mem[0819]='hd22a; mem[0820]='h070e; mem[0821]='h132d; mem[0822]='h06a0; mem[0823]='h0722; // address 0x0660
    mem[0824]='h100e; mem[0825]='h0205; mem[0826]='h0008; mem[0827]='h0878; mem[0828]='h0468; mem[0829]='h0678; mem[0830]='h0286; mem[0831]='h0047; // address 0x0670
    mem[0832]='h1106; mem[0833]='h0286; mem[0834]='h004a; mem[0835]='h1516; mem[0836]='h0226; mem[0837]='hffc9; mem[0838]='h10ec; mem[0839]='h0286; // address 0x0680
    mem[0840]='h003a; mem[0841]='h1610; mem[0842]='h04ca; mem[0843]='h0705; mem[0844]='h020c; mem[0845]='h0080; mem[0846]='h1f0f; mem[0847]='h16fb; // address 0x0690
    mem[0848]='h0605; mem[0849]='h16fc; mem[0850]='hc28a; mem[0851]='h1609; mem[0852]='h2fa0; mem[0853]='h00f2; mem[0854]='h2fa0; mem[0855]='hec02; // address 0x06a0
    mem[0856]='h0460; mem[0857]='h0142; mem[0858]='h04c0; mem[0859]='h070a; mem[0860]='h10ee; mem[0861]='hc000; mem[0862]='h1302; mem[0863]='h0460; // address 0x06b0
    mem[0864]='h0208; mem[0865]='h0460; mem[0866]='h0204; mem[0867]='h2f46; mem[0868]='h9806; mem[0869]='h00f2; mem[0870]='h16fc; mem[0871]='h10c6; // address 0x06c0
    mem[0872]='ha280; mem[0873]='hc24a; mem[0874]='h10c4; mem[0875]='ha280; mem[0876]='hce4a; mem[0877]='h10c1; mem[0878]='ha1ca; mem[0879]='h13bf; // address 0x06d0
    mem[0880]='h0200; mem[0881]='h0001; mem[0882]='h10e8; mem[0883]='h020a; mem[0884]='hec02; mem[0885]='h1003; mem[0886]='h0645; mem[0887]='h020a; // address 0x06e0
    mem[0888]='hec22; mem[0889]='h2f46; mem[0890]='hde86; mem[0891]='h0986; mem[0892]='ha1c6; mem[0893]='h0605; mem[0894]='h16fa; mem[0895]='h10af; // address 0x06f0
    mem[0896]='ha280; mem[0897]='hc38a; mem[0898]='h10ac; mem[0899]='h024a; mem[0900]='hfffe; mem[0901]='hc00a; mem[0902]='h10a8; mem[0903]='h3745; // address 0x0700
    mem[0904]='h443a; mem[0905]='h3a3a; mem[0906]='h3a32; mem[0907]='hf22d; mem[0908]='h2c30; mem[0909]='h2f47; mem[0910]='h1e00; mem[0911]='h3a3a; // address 0x0710
    mem[0912]='h3bf3; mem[0913]='h0205; mem[0914]='hfffc; mem[0915]='h1001; mem[0916]='h0705; mem[0917]='h04ca; mem[0918]='h2f46; mem[0919]='h0286; // address 0x0720
    mem[0920]='h2000; mem[0921]='h11fc; mem[0922]='h0286; mem[0923]='h5f00; mem[0924]='h15f9; mem[0925]='h0986; mem[0926]='h0288; mem[0927]='h3200; // address 0x0730
    mem[0928]='h1301; mem[0929]='ha1c6; mem[0930]='h0286; mem[0931]='h0030; mem[0932]='h1112; mem[0933]='h0286; mem[0934]='h0039; mem[0935]='h1208; // address 0x0740
    mem[0936]='h0286; mem[0937]='h0041; mem[0938]='h110c; mem[0939]='h0286; mem[0940]='h0046; mem[0941]='h1509; mem[0942]='h0226; mem[0943]='h0009; // address 0x0750
    mem[0944]='h0246; mem[0945]='h000f; mem[0946]='h0a4a; mem[0947]='ha286; mem[0948]='h0585; mem[0949]='h16e0; mem[0950]='h05cb; mem[0951]='h045b; // address 0x0760
    mem[0952]='h0203; mem[0953]='h8402; mem[0954]='h0204; mem[0955]='h05c0; mem[0956]='h0a25; mem[0957]='h1103; mem[0958]='h4008; mem[0959]='h4048; // address 0x0770
    mem[0960]='h1007; mem[0961]='h0223; mem[0962]='h1000; mem[0963]='h0224; mem[0964]='hffc0; mem[0965]='h0a82; mem[0966]='h1001; mem[0967]='h0484; // address 0x0780
    mem[0968]='h0483; mem[0969]='h1603; mem[0970]='h2fa0; mem[0971]='h00f2; mem[0972]='h2e80; mem[0973]='h8040; mem[0974]='h16f8; mem[0975]='h0459; // address 0x0790
    mem[0976]='h2fa0; mem[0977]='h00c0; mem[0978]='hc100; mem[0979]='ha101; mem[0980]='h2e84; mem[0981]='h2fa0; mem[0982]='h00c9; mem[0983]='h6001; // address 0x07a0
    mem[0984]='h2e80; mem[0985]='h0459; mem[0986]='h0560; mem[0987]='hec44; mem[0988]='h0459; mem[0989]='h04e0; mem[0990]='hec4e; mem[0991]='h04e0; // address 0x07b0
    mem[0992]='hec4c; mem[0993]='hc240; mem[0994]='h2fa0; mem[0995]='h00f2; mem[0996]='h020a; mem[0997]='h0850; mem[0998]='h0200; mem[0999]='hec52; // address 0x07c0
    mem[1000]='h0208; mem[1001]='h0006; mem[1002]='h04f0; mem[1003]='h0608; mem[1004]='h15fd; mem[1005]='h2e89; mem[1006]='h2fa0; mem[1007]='h001c; // address 0x07d0
    mem[1008]='h069a; mem[1009]='h0284; mem[1010]='h0020; mem[1011]='h1316; mem[1012]='h0284; mem[1013]='h002a; mem[1014]='h1605; mem[1015]='h069a; // address 0x07e0
    mem[1016]='h0284; mem[1017]='h000d; mem[1018]='h16fc; mem[1019]='h10e6; mem[1020]='h06a0; mem[1021]='h0bee; mem[1022]='hc807; mem[1023]='hec52; // address 0x07f0
    mem[1024]='hc809; mem[1025]='hec54; mem[1026]='hc107; mem[1027]='h06a0; mem[1028]='h0c64; mem[1029]='h1321; mem[1030]='h9807; mem[1031]='h0bf3; // address 0x0800
    mem[1032]='h1303; mem[1033]='h1004; mem[1034]='h2fa0; mem[1035]='h0021; mem[1036]='h2fa0; mem[1037]='h0021; mem[1038]='h0207; mem[1039]='h0ce3; // address 0x0810
    mem[1040]='h04c5; mem[1041]='h04c6; mem[1042]='h069a; mem[1043]='h06a0; mem[1044]='h0c34; mem[1045]='h1643; mem[1046]='h0ab4; mem[1047]='h0587; // address 0x0820
    mem[1048]='hd017; mem[1049]='h1102; mem[1050]='h1372; mem[1051]='h05c6; mem[1052]='h0a10; mem[1053]='h09e0; mem[1054]='h8005; mem[1055]='h11f7; // address 0x0830
    mem[1056]='h156c; mem[1057]='hd017; mem[1058]='h0a30; mem[1059]='h9100; mem[1060]='h16f2; mem[1061]='h0585; mem[1062]='h10eb; mem[1063]='h1065; // address 0x0840
    mem[1064]='h2f44; mem[1065]='h0284; mem[1066]='h1b00; mem[1067]='h13b6; mem[1068]='h0284; mem[1069]='h2000; mem[1070]='h1a01; mem[1071]='h2f04; // address 0x0850
    mem[1072]='h0984; mem[1073]='hc804; mem[1074]='hec60; mem[1075]='h045b; mem[1076]='h069a; mem[1077]='h0284; mem[1078]='h0027; mem[1079]='h1655; // address 0x0860
    mem[1080]='hc1c9; mem[1081]='h75d7; mem[1082]='h0588; mem[1083]='h069a; mem[1084]='h0284; mem[1085]='h0027; mem[1086]='h1358; mem[1087]='h06c4; // address 0x0870
    mem[1088]='hddc4; mem[1089]='h10f7; mem[1090]='h06a0; mem[1091]='h0b14; mem[1092]='hc806; mem[1093]='hec54; mem[1094]='h1064; mem[1095]='h070e; // address 0x0880
    mem[1096]='hc006; mem[1097]='h06a0; mem[1098]='h0b14; mem[1099]='hc809; mem[1100]='hec54; mem[1101]='h0280; mem[1102]='h0014; mem[1103]='h1605; // address 0x0890
    mem[1104]='ha189; mem[1105]='h1303; mem[1106]='h0586; mem[1107]='h8246; mem[1108]='h1a38; mem[1109]='hc246; mem[1110]='h0249; mem[1111]='hfffe; // address 0x08a0
    mem[1112]='h1052; mem[1113]='hc145; mem[1114]='h13af; mem[1115]='hd017; mem[1116]='h1130; mem[1117]='h070e; mem[1118]='h0286; mem[1119]='h0032; // address 0x08b0
    mem[1120]='h13e1; mem[1121]='h0286; mem[1122]='h009a; mem[1123]='h13d0; mem[1124]='hc026; mem[1125]='h0d76; mem[1126]='hc040; mem[1127]='h0241; // address 0x08c0
    mem[1128]='hfff0; mem[1129]='h1302; mem[1130]='hc641; mem[1131]='h05c8; mem[1132]='hc040; mem[1133]='h0241; mem[1134]='h000f; mem[1135]='hd021; // address 0x08d0
    mem[1136]='h0cd6; mem[1137]='h06c0; mem[1138]='h0260; mem[1139]='hffe0; mem[1140]='hc040; mem[1141]='h0921; mem[1142]='h0241; mem[1143]='h0006; // address 0x08e0
    mem[1144]='hc061; mem[1145]='h0cc6; mem[1146]='h1307; mem[1147]='h0284; mem[1148]='h0020; mem[1149]='h160f; mem[1150]='h04ce; mem[1151]='h020f; // address 0x08f0
    mem[1152]='h0904; mem[1153]='h0691; mem[1154]='hc040; mem[1155]='h0ad1; mem[1156]='h09c1; mem[1157]='hc061; mem[1158]='h0cc6; mem[1159]='h1309; // address 0x0900
    mem[1160]='h04c0; mem[1161]='h04ce; mem[1162]='h020f; mem[1163]='h0922; mem[1164]='h0691; mem[1165]='h2fa0; mem[1166]='h00d1; mem[1167]='h0460; // address 0x0910
    mem[1168]='h07c4; mem[1169]='h0284; mem[1170]='h000d; mem[1171]='h1307; mem[1172]='h0284; mem[1173]='h0020; mem[1174]='h16f6; mem[1175]='h069a; // address 0x0920
    mem[1176]='h0284; mem[1177]='h000d; mem[1178]='h16fc; mem[1179]='h0280; mem[1180]='h0030; mem[1181]='h135c; mem[1182]='h2f20; mem[1183]='h00f2; // address 0x0930
    mem[1184]='h2e89; mem[1185]='hc089; mem[1186]='h06a0; mem[1187]='h0c86; mem[1188]='h0204; mem[1189]='h2052; mem[1190]='hc0c3; mem[1191]='h1301; // address 0x0940
    mem[1192]='h06c4; mem[1193]='h2f04; mem[1194]='h2eb9; mem[1195]='h2fa0; mem[1196]='h00f2; mem[1197]='h0648; mem[1198]='h15f1; mem[1199]='h0200; // address 0x0950
    mem[1200]='hec56; mem[1201]='h06a0; mem[1202]='h0c9a; mem[1203]='h06a0; mem[1204]='h0c9a; mem[1205]='hc120; mem[1206]='hec52; mem[1207]='h1331; // address 0x0960
    mem[1208]='h0224; mem[1209]='h8000; mem[1210]='h06a0; mem[1211]='h0c64; mem[1212]='h1608; mem[1213]='h06a0; mem[1214]='h09d6; mem[1215]='hc390; // address 0x0970
    mem[1216]='hc403; mem[1217]='h06a0; mem[1218]='h09e6; mem[1219]='hc00e; mem[1220]='h16fa; mem[1221]='h0224; mem[1222]='h8080; mem[1223]='h06a0; // address 0x0980
    mem[1224]='h0c64; mem[1225]='h161a; mem[1226]='h06a0; mem[1227]='h09d6; mem[1228]='h04ce; mem[1229]='h0580; mem[1230]='hd390; mem[1231]='hc083; // address 0x0990
    mem[1232]='h6080; mem[1233]='h0602; mem[1234]='h0a72; mem[1235]='h1907; mem[1236]='h0600; mem[1237]='h2e80; mem[1238]='h2fa0; mem[1239]='h00d1; // address 0x09a0
    mem[1240]='h2fa0; mem[1241]='h00f2; mem[1242]='h1004; mem[1243]='hd402; mem[1244]='h0600; mem[1245]='h06a0; mem[1246]='h09e6; mem[1247]='h087e; // address 0x09b0
    mem[1248]='h05ce; mem[1249]='h1302; mem[1250]='ha00e; mem[1251]='h10e8; mem[1252]='h0200; mem[1253]='hec52; mem[1254]='h04c4; mem[1255]='h06a0; // address 0x09c0
    mem[1256]='h0c9c; mem[1257]='h0460; mem[1258]='h07c8; mem[1259]='hc012; mem[1260]='h04e2; mem[1261]='hfffe; mem[1262]='h0620; mem[1263]='hec4c; // address 0x09d0
    mem[1264]='hc0e0; mem[1265]='hec54; mem[1266]='h045b; mem[1267]='h2e80; mem[1268]='h2f20; mem[1269]='h0a05; mem[1270]='h2e90; mem[1271]='h2fa0; // address 0x09e0
    mem[1272]='h00f2; mem[1273]='h045b; mem[1274]='h2fa0; mem[1275]='h001f; mem[1276]='h2ea0; mem[1277]='hec4c; mem[1278]='h0460; mem[1279]='h0142; // address 0x09f0
    mem[1280]='h069a; mem[1281]='h0284; mem[1282]='h002a; mem[1283]='h131a; mem[1284]='h0284; mem[1285]='h0040; mem[1286]='h1622; mem[1287]='h06a0; // address 0x0a00
    mem[1288]='h0b14; mem[1289]='hc088; mem[1290]='ha089; mem[1291]='hc486; mem[1292]='h05c8; mem[1293]='h0206; mem[1294]='h0020; mem[1295]='h0284; // address 0x0a10
    mem[1296]='h0028; mem[1297]='h1608; mem[1298]='h06a0; mem[1299]='h0ad0; mem[1300]='h0266; mem[1301]='h0020; mem[1302]='h0284; mem[1303]='h0029; // address 0x0a20
    mem[1304]='h1649; mem[1305]='h069a; mem[1306]='hc000; mem[1307]='h1601; mem[1308]='h0a66; mem[1309]='h1040; mem[1310]='h06a0; mem[1311]='h0ad0; // address 0x0a30
    mem[1312]='h0266; mem[1313]='h0010; mem[1314]='h0284; mem[1315]='h002b; mem[1316]='h1603; mem[1317]='h069a; mem[1318]='h0266; mem[1319]='h0030; // address 0x0a40
    mem[1320]='h10f1; mem[1321]='h020e; mem[1322]='h0a34; mem[1323]='hc80e; mem[1324]='hec5e; mem[1325]='h0460; mem[1326]='h0ad6; mem[1327]='h06a0; // address 0x0a50
    mem[1328]='h0ad0; mem[1329]='h0a46; mem[1330]='h102b; mem[1331]='hc006; mem[1332]='h0280; mem[1333]='h0030; mem[1334]='h1604; mem[1335]='h0284; // address 0x0a60
    mem[1336]='h000d; mem[1337]='h1312; mem[1338]='h070e; mem[1339]='h06a0; mem[1340]='h0b14; mem[1341]='h0280; mem[1342]='h0030; mem[1343]='h130b; // address 0x0a70
    mem[1344]='hc089; mem[1345]='ha088; mem[1346]='hc486; mem[1347]='h05c8; mem[1348]='h0280; mem[1349]='h0026; mem[1350]='h1605; mem[1351]='h070e; // address 0x0a80
    mem[1352]='h0284; mem[1353]='h002c; mem[1354]='h13f0; mem[1355]='hc386; mem[1356]='h045f; mem[1357]='h06a0; mem[1358]='h0ad0; mem[1359]='h10ca; // address 0x0a90
    mem[1360]='h06a0; mem[1361]='h0b14; mem[1362]='hc089; mem[1363]='h05c2; mem[1364]='h6182; mem[1365]='h0816; mem[1366]='h0286; mem[1367]='h007f; // address 0x0aa0
    mem[1368]='h1507; mem[1369]='h0286; mem[1370]='hff80; mem[1371]='h1104; mem[1372]='h0246; mem[1373]='h00ff; mem[1374]='he646; mem[1375]='h045f; // address 0x0ab0
    mem[1376]='h2fa0; mem[1377]='h00d6; mem[1378]='h0460; mem[1379]='h091a; mem[1380]='h070e; mem[1381]='h06a0; mem[1382]='h0b14; mem[1383]='h10ee; // address 0x0ac0
    mem[1384]='hc80b; mem[1385]='hec5e; mem[1386]='h069a; mem[1387]='h020c; mem[1388]='h0b04; mem[1389]='h0284; mem[1390]='h0052; mem[1391]='h130c; // address 0x0ad0
    mem[1392]='h0284; mem[1393]='h003a; mem[1394]='h110a; mem[1395]='h0284; mem[1396]='h003e; mem[1397]='h1309; mem[1398]='h020e; mem[1399]='hfffe; // address 0x0ae0
    mem[1400]='h020d; mem[1401]='h0b04; mem[1402]='h0460; mem[1403]='h0b18; mem[1404]='h069a; mem[1405]='h0460; mem[1406]='h0c2a; mem[1407]='h069a; // address 0x0af0
    mem[1408]='h0460; mem[1409]='h0c0c; mem[1410]='hc145; mem[1411]='h11de; mem[1412]='h0286; mem[1413]='h0010; mem[1414]='h14db; mem[1415]='hc2e0; // address 0x0b00
    mem[1416]='hec5e; mem[1417]='h045b; mem[1418]='hc34b; mem[1419]='h069a; mem[1420]='h04e0; mem[1421]='hec50; mem[1422]='h0284; mem[1423]='h0027; // address 0x0b10
    mem[1424]='h1307; mem[1425]='h0284; mem[1426]='h002d; mem[1427]='h1610; mem[1428]='h054d; mem[1429]='h05ce; mem[1430]='h069a; mem[1431]='h1011; // address 0x0b20
    mem[1432]='h04c6; mem[1433]='h04ce; mem[1434]='h069a; mem[1435]='h0284; mem[1436]='h0027; mem[1437]='h1304; mem[1438]='h06c6; mem[1439]='hd106; // address 0x0b30
    mem[1440]='hc184; mem[1441]='h10f8; mem[1442]='h069a; mem[1443]='h1043; mem[1444]='h0284; mem[1445]='h002b; mem[1446]='h13ee; mem[1447]='hc38e; // address 0x0b40
    mem[1448]='h154b; mem[1449]='h0284; mem[1450]='h0024; mem[1451]='h1603; mem[1452]='hc189; mem[1453]='h069a; mem[1454]='h1037; mem[1455]='h0284; // address 0x0b50
    mem[1456]='h003e; mem[1457]='h1604; mem[1458]='h069a; mem[1459]='h06a0; mem[1460]='h0c0a; mem[1461]='h1030; mem[1462]='h06a0; mem[1463]='h0c34; // address 0x0b60
    mem[1464]='h11a9; mem[1465]='h1325; mem[1466]='h06a0; mem[1467]='h0c28; mem[1468]='h1029; mem[1469]='hc38e; mem[1470]='h16a3; mem[1471]='hc059; // address 0x0b70
    mem[1472]='h04c2; mem[1473]='h06a0; mem[1474]='h0c86; mem[1475]='hc4c9; mem[1476]='h0241; mem[1477]='hf000; mem[1478]='h0281; mem[1479]='h1000; // address 0x0b80
    mem[1480]='h1611; mem[1481]='h0264; mem[1482]='h0080; mem[1483]='hc189; mem[1484]='h0643; mem[1485]='hc4c4; mem[1486]='h8820; mem[1487]='hec56; // address 0x0b90
    mem[1488]='hec5a; mem[1489]='h1603; mem[1490]='hc1a0; mem[1491]='hec58; mem[1492]='h1012; mem[1493]='h06a0; mem[1494]='h0c64; mem[1495]='h1601; // address 0x0ba0
    mem[1496]='hc192; mem[1497]='h100d; mem[1498]='ha4c8; mem[1499]='h0264; mem[1500]='h8000; mem[1501]='h04c6; mem[1502]='h10ed; mem[1503]='h06a0; // address 0x0bb0
    mem[1504]='h0bee; mem[1505]='hc107; mem[1506]='h06a0; mem[1507]='h0c64; mem[1508]='h16d8; mem[1509]='hc192; mem[1510]='h05ce; mem[1511]='hc120; // address 0x0bc0
    mem[1512]='hec60; mem[1513]='hc34d; mem[1514]='h1502; mem[1515]='h0506; mem[1516]='h054d; mem[1517]='hc145; mem[1518]='h1194; mem[1519]='hc38e; // address 0x0bd0
    mem[1520]='h1305; mem[1521]='ha806; mem[1522]='hec50; mem[1523]='h109d; mem[1524]='hc1a0; mem[1525]='hec50; mem[1526]='h045d; mem[1527]='hc30b; // address 0x0be0
    mem[1528]='h0207; mem[1529]='h0031; mem[1530]='h06a0; mem[1531]='h0c34; mem[1532]='h111c; mem[1533]='h1303; mem[1534]='h0a87; mem[1535]='h1919; // address 0x0bf0
    mem[1536]='h1001; mem[1537]='h0a87; mem[1538]='ha1c4; mem[1539]='h069a; mem[1540]='h10f5; mem[1541]='hc30b; mem[1542]='h0202; mem[1543]='h0010; // address 0x0c00
    mem[1544]='h04c6; mem[1545]='h0705; mem[1546]='h06a0; mem[1547]='h0c34; mem[1548]='h110c; mem[1549]='h8083; mem[1550]='h1409; mem[1551]='hc146; // address 0x0c10
    mem[1552]='h3942; mem[1553]='ha183; mem[1554]='h069a; mem[1555]='h10f6; mem[1556]='hc30b; mem[1557]='h0202; mem[1558]='h000a; mem[1559]='h10f0; // address 0x0c20
    mem[1560]='h0705; mem[1561]='h045c; mem[1562]='h0701; mem[1563]='hc0c4; mem[1564]='h0284; mem[1565]='h0024; mem[1566]='h1306; mem[1567]='h0223; // address 0x0c30
    mem[1568]='hffd0; mem[1569]='h170e; mem[1570]='h0283; mem[1571]='h0009; mem[1572]='h1502; mem[1573]='h0501; mem[1574]='h045b; mem[1575]='h0223; // address 0x0c40
    mem[1576]='hfff9; mem[1577]='h0283; mem[1578]='h000a; mem[1579]='h1a04; mem[1580]='h0283; mem[1581]='h0023; mem[1582]='h1b01; mem[1583]='h04c1; // address 0x0c50
    mem[1584]='hc041; mem[1585]='h045b; mem[1586]='h0703; mem[1587]='hc060; mem[1588]='hec4e; mem[1589]='h130b; mem[1590]='h0a21; mem[1591]='h0202; // address 0x0c60
    mem[1592]='hec62; mem[1593]='ha042; mem[1594]='h04c3; mem[1595]='h05c2; mem[1596]='h8c84; mem[1597]='h1303; mem[1598]='h8042; mem[1599]='h1afb; // address 0x0c70
    mem[1600]='h0583; mem[1601]='hc0c3; mem[1602]='h045b; mem[1603]='h0203; mem[1604]='hec58; mem[1605]='h84c2; mem[1606]='h1305; mem[1607]='h0203; // address 0x0c80
    mem[1608]='hec5c; mem[1609]='h84c2; mem[1610]='h1301; mem[1611]='h04c3; mem[1612]='h045b; mem[1613]='hc110; mem[1614]='hc30b; mem[1615]='h06a0; // address 0x0c90
    mem[1616]='h0c64; mem[1617]='h130d; mem[1618]='hc104; mem[1619]='h1304; mem[1620]='h04c4; mem[1621]='h05a0; mem[1622]='hec4c; mem[1623]='h10f7; // address 0x0ca0
    mem[1624]='h05a0; mem[1625]='hec4e; mem[1626]='hc0a0; mem[1627]='hec4e; mem[1628]='h0a22; mem[1629]='h0222; mem[1630]='hec62; mem[1631]='h0642; // address 0x0cb0
    mem[1632]='hccb0; mem[1633]='hc4b0; mem[1634]='h045c; mem[1635]='h0000; mem[1636]='h0a00; mem[1637]='h0a9a; mem[1638]='h0a66; mem[1639]='h0a5e; // address 0x0cc0
    mem[1640]='h0aa0; mem[1641]='h0ac8; mem[1642]='h088e; mem[1643]='h0905; mem[1644]='h0a0a; mem[1645]='h1408; mem[1646]='h0013; mem[1647]='h0a06; // address 0x0cd0
    mem[1648]='h0310; mem[1649]='h0307; mem[1650]='h0122; mem[1651]='h5329; mem[1652]='haec4; mem[1653]='h69af; mem[1654]='hd267; mem[1655]='h022c; // address 0x0ce0
    mem[1656]='hd770; mem[1657]='hb353; mem[1658]='h0322; mem[1659]='h29ab; mem[1660]='hcf6e; mem[1661]='h66ac; mem[1662]='h52af; mem[1663]='h43ba; // address 0x0cf0
    mem[1664]='h4384; mem[1665]='ha1d4; mem[1666]='h61a5; mem[1667]='h4374; mem[1668]='ha956; mem[1669]='h7385; mem[1670]='hae44; mem[1671]='hb155; // address 0x0d00
    mem[1672]='h89a4; mem[1673]='hcc65; mem[1674]='hae43; mem[1675]='h7456; mem[1676]='h8aa5; mem[1677]='h51a7; mem[1678]='h5428; mem[1679]='h452c; // address 0x0d10
    mem[1680]='h4554; mem[1681]='had50; mem[1682]='hae43; mem[1683]='h454f; mem[1684]='haf43; mem[1685]='h508c; mem[1686]='ha4c3; mem[1687]='h7229; // address 0x0d20
    mem[1688]='hcd69; mem[1689]='hb2c5; mem[1690]='h78b3; mem[1691]='h54b7; mem[1692]='h5069; mem[1693]='h8daf; mem[1694]='h5662; mem[1695]='hb059; // address 0x0d30
    mem[1696]='h738e; mem[1697]='ha547; mem[1698]='haf50; mem[1699]='h8fb2; mem[1700]='h4992; mem[1701]='hb3c5; mem[1702]='h74b4; mem[1703]='hd770; // address 0x0d40
    mem[1704]='h1322; mem[1705]='h4f5a; mem[1706]='ha5d4; mem[1707]='h6fac; mem[1708]='h41af; mem[1709]='h4362; mem[1710]='hb241; mem[1711]='h434c; // address 0x0d50
    mem[1712]='hb4c3; mem[1713]='h72d3; mem[1714]='h74d7; mem[1715]='h70b7; mem[1716]='hd062; mem[1717]='hba43; mem[1718]='h6294; mem[1719]='h22a5; // address 0x0d60
    mem[1720]='hd874; mem[1721]='h18af; mem[1722]='h5052; mem[1723]='h0000; mem[1724]='ha000; mem[1725]='hb000; mem[1726]='h0745; mem[1727]='h0227; // address 0x0d70
    mem[1728]='h0247; mem[1729]='h000d; mem[1730]='h0445; mem[1731]='h0685; mem[1732]='h0405; mem[1733]='h000d; mem[1734]='h8000; mem[1735]='h9000; // address 0x0d80
    mem[1736]='h0287; mem[1737]='h03a6; mem[1738]='h03c6; mem[1739]='h04c5; mem[1740]='h2002; mem[1741]='h2402; mem[1742]='h000a; mem[1743]='h0605; // address 0x0d90
    mem[1744]='h0645; mem[1745]='h3c08; mem[1746]='h0185; mem[1747]='h000c; mem[1748]='h0006; mem[1749]='h0346; mem[1750]='h0585; mem[1751]='h05c5; // address 0x0da0
    mem[1752]='h0545; mem[1753]='h1301; mem[1754]='h1501; mem[1755]='h1b01; mem[1756]='h1401; mem[1757]='h1a01; mem[1758]='h1201; mem[1759]='h1101; // address 0x0db0
    mem[1760]='h1001; mem[1761]='h1701; mem[1762]='h1601; mem[1763]='h1901; mem[1764]='h1801; mem[1765]='h1c01; mem[1766]='h3003; mem[1767]='h0207; // address 0x0dc0
    mem[1768]='h030a; mem[1769]='h03e6; mem[1770]='h008b; mem[1771]='h009b; mem[1772]='h02ea; mem[1773]='hc000; mem[1774]='hd000; mem[1775]='h3808; // address 0x0dd0
    mem[1776]='h01c5; mem[1777]='h0505; mem[1778]='h1006; mem[1779]='h0267; mem[1780]='h0366; mem[1781]='h0386; mem[1782]='h6000; mem[1783]='h7000; // address 0x0de0
    mem[1784]='h1d09; mem[1785]='h1e09; mem[1786]='h0705; mem[1787]='h0a04; mem[1788]='he000; mem[1789]='hf000; mem[1790]='h0804; mem[1791]='h0b04; // address 0x0df0
    mem[1792]='h0904; mem[1793]='h3403; mem[1794]='h02cb; mem[1795]='h02ab; mem[1796]='h06c5; mem[1797]='h4000; mem[1798]='h5000; mem[1799]='h1f09; // address 0x0e00
    mem[1800]='h0006; mem[1801]='h0485; mem[1802]='h2c08; mem[1803]='h2802; mem[1804]='h0000; mem[1805]='h02e0; mem[1806]='hec00; mem[1807]='h0203; // address 0x0e10
    mem[1808]='hec4c; mem[1809]='h0205; mem[1810]='hed00; mem[1811]='h0206; mem[1812]='heffe; mem[1813]='hccc5; mem[1814]='hccc6; mem[1815]='hccc5; // address 0x0e20
    mem[1816]='h04c5; mem[1817]='h04d3; mem[1818]='h0209; mem[1819]='hec2e; mem[1820]='hc820; mem[1821]='hec44; mem[1822]='hec54; mem[1823]='h020c; // address 0x0e30
    mem[1824]='h0400; mem[1825]='h1d1f; mem[1826]='h3220; mem[1827]='h013b; mem[1828]='h1e0d; mem[1829]='h3320; mem[1830]='h0096; mem[1831]='h1d10; // address 0x0e40
    mem[1832]='h020c; mem[1833]='h0000; mem[1834]='h1d0e; mem[1835]='h3220; mem[1836]='h013b; mem[1837]='h04c1; mem[1838]='h04c2; mem[1839]='hc660; // address 0x0e50
    mem[1840]='h013e; mem[1841]='h2fa0; mem[1842]='h00e3; mem[1843]='h05e0; mem[1844]='hec44; mem[1845]='h020c; mem[1846]='h0000; mem[1847]='h1f15; // address 0x0e60
    mem[1848]='h1334; mem[1849]='h020c; mem[1850]='h0400; mem[1851]='h1f15; mem[1852]='h1303; mem[1853]='hc041; mem[1854]='h162c; mem[1855]='h10f5; // address 0x0e70
    mem[1856]='hc660; mem[1857]='h0140; mem[1858]='hc082; mem[1859]='h1625; mem[1860]='h2f4a; mem[1861]='h028a; mem[1862]='h0000; mem[1863]='h13ed; // address 0x0e80
    mem[1864]='h028a; mem[1865]='h7f00; mem[1866]='h13ea; mem[1867]='h028a; mem[1868]='h1000; mem[1869]='h160d; mem[1870]='h2f4a; mem[1871]='h028a; // address 0x0e90
    mem[1872]='h0000; mem[1873]='h13fc; mem[1874]='h028a; mem[1875]='h3700; mem[1876]='h130e; mem[1877]='h028a; mem[1878]='h3c00; mem[1879]='h16dd; // address 0x0ea0
    mem[1880]='h2f20; mem[1881]='h013c; mem[1882]='h10da; mem[1883]='h028a; mem[1884]='h1200; mem[1885]='h1602; mem[1886]='h0460; mem[1887]='h1070; // address 0x0eb0
    mem[1888]='h028a; mem[1889]='h1100; mem[1890]='h1602; mem[1891]='h0460; mem[1892]='h0fa0; mem[1893]='hc660; mem[1894]='h013e; mem[1895]='h2f0a; // address 0x0ec0
    mem[1896]='h10cc; mem[1897]='h0460; mem[1898]='h107c; mem[1899]='h0460; mem[1900]='h0fc8; mem[1901]='hc660; mem[1902]='h013e; mem[1903]='h2f4a; // address 0x0ed0
    mem[1904]='h028a; mem[1905]='h1a00; mem[1906]='h1605; mem[1907]='hc820; mem[1908]='hec54; mem[1909]='hec44; mem[1910]='h0460; mem[1911]='h0142; // address 0x0ee0
    mem[1912]='h028a; mem[1913]='h0300; mem[1914]='h1310; mem[1915]='h028a; mem[1916]='h1200; mem[1917]='h13e0; mem[1918]='h028a; mem[1919]='h1400; // address 0x0ef0
    mem[1920]='h1602; mem[1921]='h0460; mem[1922]='h10fe; mem[1923]='hc041; mem[1924]='h16e6; mem[1925]='hc082; mem[1926]='h16e2; mem[1927]='hc660; // address 0x0f00
    mem[1928]='h0140; mem[1929]='h2f0a; mem[1930]='h10aa; mem[1931]='hc660; mem[1932]='h013e; mem[1933]='hc820; mem[1934]='hec54; mem[1935]='hec44; // address 0x0f10
    mem[1936]='h2fa0; mem[1937]='h00d8; mem[1938]='h2eca; mem[1939]='h2fa0; mem[1940]='h00de; mem[1941]='h06a0; mem[1942]='h0f42; mem[1943]='h5500; // address 0x0f20
    mem[1944]='h0f7e; mem[1945]='h4400; mem[1946]='h0f94; mem[1947]='h5400; mem[1948]='h0f5a; mem[1949]='h5100; mem[1950]='h0e5a; mem[1951]='h0000; // address 0x0f30
    mem[1952]='h05cb; mem[1953]='hc01b; mem[1954]='h1304; mem[1955]='h82bb; mem[1956]='h16fb; mem[1957]='hc2db; mem[1958]='h045b; mem[1959]='h2fa0; // address 0x0f40
    mem[1960]='h00f5; mem[1961]='h10e1; mem[1962]='h2fa0; mem[1963]='h00ff; mem[1964]='h10de; mem[1965]='h2e4a; mem[1966]='h0f16; mem[1967]='h0f54; // address 0x0f50
    mem[1968]='h0a2a; mem[1969]='h064a; mem[1970]='h12f7; mem[1971]='h028a; mem[1972]='h0023; mem[1973]='h14f4; mem[1974]='h020c; mem[1975]='h0400; // address 0x0f60
    mem[1976]='h1d0b; mem[1977]='h1d0c; mem[1978]='h332a; mem[1979]='h0084; mem[1980]='h1e0b; mem[1981]='h1e0c; mem[1982]='h10cc; mem[1983]='h2e4a; // address 0x0f70
    mem[1984]='h0f88; mem[1985]='h0f54; mem[1986]='hc80a; mem[1987]='hec50; mem[1988]='h2e4a; mem[1989]='h0f16; mem[1990]='h0f54; mem[1991]='hc80a; // address 0x0f80
    mem[1992]='hec4e; mem[1993]='h10c1; mem[1994]='h2e4a; mem[1995]='h0f16; mem[1996]='h0f54; mem[1997]='hc80a; mem[1998]='hec4c; mem[1999]='h10bb; // address 0x0f90
    mem[2000]='h0701; mem[2001]='hc1e0; mem[2002]='hec52; mem[2003]='h112d; mem[2004]='h1533; mem[2005]='hc1e0; mem[2006]='hec50; mem[2007]='h8807; // address 0x0fa0
    mem[2008]='hec4e; mem[2009]='h1b37; mem[2010]='hc660; mem[2011]='h0140; mem[2012]='h04c5; mem[2013]='h04c3; mem[2014]='h2fa0; mem[2015]='h0137; // address 0x0fb0
    mem[2016]='hc287; mem[2017]='h06a0; mem[2018]='h1042; mem[2019]='h3900; mem[2020]='hc297; mem[2021]='h06a0; mem[2022]='h1042; mem[2023]='h4200; // address 0x0fc0
    mem[2024]='h8807; mem[2025]='hec4e; mem[2026]='h1a03; mem[2027]='h0720; mem[2028]='hec52; mem[2029]='h1004; mem[2030]='h05c7; mem[2031]='h0283; // address 0x0fd0
    mem[2032]='h003c; mem[2033]='h111d; mem[2034]='h0225; mem[2035]='h0037; mem[2036]='hc285; mem[2037]='h050a; mem[2038]='h06a0; mem[2039]='h1042; // address 0x0fe0
    mem[2040]='h3700; mem[2041]='hc807; mem[2042]='hec50; mem[2043]='h2fa0; mem[2044]='h0128; mem[2045]='hc160; mem[2046]='hec54; mem[2047]='h110e; // address 0x0ff0
    mem[2048]='h10cf; mem[2049]='h2fa0; mem[2050]='h0137; mem[2051]='h2fa0; mem[2052]='h00e0; mem[2053]='h05e0; mem[2054]='hec52; mem[2055]='h10f5; // address 0x1000
    mem[2056]='h2fa0; mem[2057]='h0137; mem[2058]='h2fa0; mem[2059]='h0131; mem[2060]='h04e0; mem[2061]='hec52; mem[2062]='h04c1; mem[2063]='h0460; // address 0x1010
    mem[2064]='h0e6a; mem[2065]='h2fa0; mem[2066]='h0137; mem[2067]='h2fa0; mem[2068]='h0131; mem[2069]='hc660; mem[2070]='h013e; mem[2071]='hc820; // address 0x1020
    mem[2072]='hec54; mem[2073]='hec44; mem[2074]='h2fa0; mem[2075]='h011f; mem[2076]='h05e0; mem[2077]='hec44; mem[2078]='h0720; mem[2079]='hec4c; // address 0x1030
    mem[2080]='h10eb; mem[2081]='hc03b; mem[2082]='h2f00; mem[2083]='h0980; mem[2084]='ha140; mem[2085]='h2e8a; mem[2086]='h0223; mem[2087]='h0005; // address 0x1040
    mem[2088]='h0200; mem[2089]='h0004; mem[2090]='h0b4a; mem[2091]='hc18a; mem[2092]='h09c6; mem[2093]='ha146; mem[2094]='h0225; mem[2095]='h0030; // address 0x1050
    mem[2096]='h0286; mem[2097]='h000a; mem[2098]='h1a02; mem[2099]='h0225; mem[2100]='h0007; mem[2101]='h0600; mem[2102]='h16f3; mem[2103]='h045b; // address 0x1060
    mem[2104]='h0702; mem[2105]='hc660; mem[2106]='h0140; mem[2107]='hc020; mem[2108]='hec4c; mem[2109]='h04c7; mem[2110]='h2f46; mem[2111]='h0286; // address 0x1070
    mem[2112]='h1400; mem[2113]='h133d; mem[2114]='hc220; mem[2115]='hec52; mem[2116]='h1657; mem[2117]='h0286; mem[2118]='h2000; mem[2119]='h11f6; // address 0x1080
    mem[2120]='h0286; mem[2121]='h5f00; mem[2122]='h15f3; mem[2123]='h0705; mem[2124]='h04ca; mem[2125]='h06a0; mem[2126]='h073a; mem[2127]='h100b; // address 0x1090
    mem[2128]='hd22a; mem[2129]='h1152; mem[2130]='h1332; mem[2131]='h06a0; mem[2132]='h0722; mem[2133]='h100e; mem[2134]='h0205; mem[2135]='h0008; // address 0x10a0
    mem[2136]='h0878; mem[2137]='h0468; mem[2138]='h10b2; mem[2139]='h0286; mem[2140]='h0047; mem[2141]='h1106; mem[2142]='h0286; mem[2143]='h004a; // address 0x10b0
    mem[2144]='h1522; mem[2145]='h0226; mem[2146]='hffc9; mem[2147]='h10ec; mem[2148]='h0286; mem[2149]='h003a; mem[2150]='h161c; mem[2151]='h103e; // address 0x10c0
    mem[2152]='h020c; mem[2153]='h0400; mem[2154]='h04c5; mem[2155]='h1f0f; mem[2156]='h16fd; mem[2157]='h0605; mem[2158]='h16fc; mem[2159]='hc660; // address 0x10d0
    mem[2160]='h013e; mem[2161]='hc820; mem[2162]='hec54; mem[2163]='hec44; mem[2164]='h0720; mem[2165]='hec4c; mem[2166]='hc000; mem[2167]='h1303; // address 0x10e0
    mem[2168]='h2fa0; mem[2169]='h010a; mem[2170]='h1002; mem[2171]='h2fa0; mem[2172]='h0115; mem[2173]='h05e0; mem[2174]='hec44; mem[2175]='h04c2; // address 0x10f0
    mem[2176]='h04e0; mem[2177]='hec52; mem[2178]='h1021; mem[2179]='h04c0; mem[2180]='h10e3; mem[2181]='h2f46; mem[2182]='h9806; mem[2183]='h00f2; // address 0x1100
    mem[2184]='h16fc; mem[2185]='h04c7; mem[2186]='h1019; mem[2187]='ha1ca; mem[2188]='h1317; mem[2189]='h0700; mem[2190]='h10d9; mem[2191]='ha280; // address 0x1110
    mem[2192]='hc0ca; mem[2193]='h1012; mem[2194]='ha280; mem[2195]='hccca; mem[2196]='h100f; mem[2197]='h0645; mem[2198]='h2f46; mem[2199]='h0986; // address 0x1120
    mem[2200]='h13fd; mem[2201]='ha1c6; mem[2202]='h0605; mem[2203]='h16fa; mem[2204]='h1007; mem[2205]='ha280; mem[2206]='hc80a; mem[2207]='hec1c; // address 0x1130
    mem[2208]='h1003; mem[2209]='h024a; mem[2210]='hfffe; mem[2211]='hc00a; mem[2212]='h0460; mem[2213]='h0e6a; mem[2214]='h0720; mem[2215]='hec52; // address 0x1140
    mem[2216]='h10fb; mem[2217]='h3d45; mem[2218]='h443c; mem[2219]='h3c3c; mem[2220]='h3c32; mem[2221]='he437; mem[2222]='h363a; mem[2223]='h3948; // address 0x1150
    mem[2224]='h2a00; mem[2225]='h3c3c; mem[2226]='h3d8b; mem[2227]='hc141; mem[2228]='h0208; mem[2229]='h12d8; mem[2230]='h0209; mem[2231]='h12ba; // address 0x1160
    mem[2232]='h0207; mem[2233]='h12a6; mem[2234]='h2fa0; mem[2235]='h00f2; mem[2236]='h0206; mem[2237]='h202c; mem[2238]='hc050; mem[2239]='h2e80; // address 0x1170
    mem[2240]='h2f06; mem[2241]='h2e81; mem[2242]='h2f06; mem[2243]='h04c3; mem[2244]='hc050; mem[2245]='h0241; mem[2246]='hfff0; mem[2247]='hc2a3; // address 0x1180
    mem[2248]='h13b4; mem[2249]='hc08a; mem[2250]='h1329; mem[2251]='h024a; mem[2252]='hfff0; mem[2253]='h8281; mem[2254]='h1402; mem[2255]='h0643; // address 0x1190
    mem[2256]='h10f6; mem[2257]='hc050; mem[2258]='h0a13; mem[2259]='h0223; mem[2260]='h14d6; mem[2261]='h604a; mem[2262]='h0242; mem[2263]='h000f; // address 0x11a0
    mem[2264]='hd0a2; mem[2265]='h11ba; mem[2266]='h0972; mem[2267]='h0462; mem[2268]='h11ba; mem[2269]='h060c; mem[2270]='h061f; mem[2271]='h232b; // address 0x11b0
    mem[2272]='h3337; mem[2273]='h063f; mem[2274]='h4145; mem[2275]='h0697; mem[2276]='h0698; mem[2277]='h2f06; mem[2278]='h0961; mem[2279]='h0698; // address 0x11c0
    mem[2280]='h103d; mem[2281]='hc041; mem[2282]='h1603; mem[2283]='h0203; mem[2284]='h14da; mem[2285]='h1024; mem[2286]='h06c1; mem[2287]='h0871; // address 0x11d0
    mem[2288]='h05c1; mem[2289]='ha040; mem[2290]='h0697; mem[2291]='h1004; mem[2292]='hc050; mem[2293]='h0203; mem[2294]='h14de; mem[2295]='h0697; // address 0x11e0
    mem[2296]='h2f20; mem[2297]='h14f5; mem[2298]='h2e81; mem[2299]='h102a; mem[2300]='h0697; mem[2301]='h0698; mem[2302]='hc209; mem[2303]='h10e5; // address 0x11f0
    mem[2304]='hd041; mem[2305]='h16f2; mem[2306]='h0b41; mem[2307]='hd081; mem[2308]='h0a61; mem[2309]='h09c2; mem[2310]='ha042; mem[2311]='h10f4; // address 0x1200
    mem[2312]='h8810; mem[2313]='h1320; mem[2314]='h1603; mem[2315]='h0203; mem[2316]='h14ee; mem[2317]='h1004; mem[2318]='h0697; mem[2319]='h10d7; // address 0x1210
    mem[2320]='hc041; mem[2321]='h16e2; mem[2322]='h0697; mem[2323]='h1012; mem[2324]='h0ac1; mem[2325]='h18de; mem[2326]='h09c1; mem[2327]='h0697; // address 0x1220
    mem[2328]='h0698; mem[2329]='h2f06; mem[2330]='hc070; mem[2331]='h10dc; mem[2332]='h0697; mem[2333]='h1019; mem[2334]='hc041; mem[2335]='h16d4; // address 0x1230
    mem[2336]='h0697; mem[2337]='h10f8; mem[2338]='h0ac1; mem[2339]='h18d0; mem[2340]='h09c1; mem[2341]='h10e2; mem[2342]='hc145; mem[2343]='h1603; // address 0x1240
    mem[2344]='hc740; mem[2345]='h0460; mem[2346]='h0142; mem[2347]='hc320; mem[2348]='h013e; mem[2349]='h1f15; mem[2350]='h1604; mem[2351]='h2f42; // address 0x1250
    mem[2352]='h0282; mem[2353]='h2f00; mem[2354]='h13f5; mem[2355]='h8140; mem[2356]='h1bf3; mem[2357]='h0460; mem[2358]='h1168; mem[2359]='h0203; // address 0x1260
    mem[2360]='h2d31; mem[2361]='h06c1; mem[2362]='h0881; mem[2363]='h1315; mem[2364]='h1502; mem[2365]='h2f03; mem[2366]='h0501; mem[2367]='h0281; // address 0x1270
    mem[2368]='h0064; mem[2369]='h1104; mem[2370]='h0a83; mem[2371]='h2f03; mem[2372]='h0221; mem[2373]='hff9c; mem[2374]='h0204; mem[2375]='h000a; // address 0x1280
    mem[2376]='hc081; mem[2377]='h04c1; mem[2378]='h3c44; mem[2379]='h0a83; mem[2380]='h1302; mem[2381]='hc041; mem[2382]='h1301; mem[2383]='h0699; // address 0x1290
    mem[2384]='hc042; mem[2385]='h0699; mem[2386]='h10d3; mem[2387]='h0202; mem[2388]='h0004; mem[2389]='h2f13; mem[2390]='h0583; mem[2391]='h0602; // address 0x12a0
    mem[2392]='h16fc; mem[2393]='h2f06; mem[2394]='h06c6; mem[2395]='h05c0; mem[2396]='h045b; mem[2397]='hc0c1; mem[2398]='h0ac3; mem[2399]='h0943; // address 0x12b0
    mem[2400]='h0283; mem[2401]='h0900; mem[2402]='h1203; mem[2403]='h06c3; mem[2404]='h0223; mem[2405]='h0126; mem[2406]='h0223; mem[2407]='h3000; // address 0x12c0
    mem[2408]='h2f03; mem[2409]='h0a83; mem[2410]='h16fd; mem[2411]='h045b; mem[2412]='h0204; mem[2413]='h2a52; mem[2414]='hc081; mem[2415]='h0aa2; // address 0x12d0
    mem[2416]='h09e2; mem[2417]='h1603; mem[2418]='h06c4; mem[2419]='h2f04; mem[2420]='h10e8; mem[2421]='h0602; mem[2422]='h1602; mem[2423]='h2f04; // address 0x12e0
    mem[2424]='h10f9; mem[2425]='h0602; mem[2426]='h1610; mem[2427]='h2fa0; mem[2428]='h14f4; mem[2429]='h2eb0; mem[2430]='hc081; mem[2431]='h0ac2; // address 0x12f0
    mem[2432]='h13ea; mem[2433]='h0202; mem[2434]='h2829; mem[2435]='h2f02; mem[2436]='h06c4; mem[2437]='h2f04; mem[2438]='hc30b; mem[2439]='h0699; // address 0x1300
    mem[2440]='h06c2; mem[2441]='h2f02; mem[2442]='h045c; mem[2443]='h2fa0; mem[2444]='h14f7; mem[2445]='h0202; mem[2446]='h002b; mem[2447]='h10f6; // address 0x1310
    mem[2448]='h045b; mem[2449]='h0000; mem[2450]='h008b; mem[2451]='h009b; mem[2452]='h0185; mem[2453]='h01c5; mem[2454]='h0207; mem[2455]='h0227; // address 0x1320
    mem[2456]='h0247; mem[2457]='h0267; mem[2458]='h0287; mem[2459]='h02ab; mem[2460]='h02cb; mem[2461]='h02ea; mem[2462]='h030a; mem[2463]='h0346; // address 0x1330
    mem[2464]='h0366; mem[2465]='h0386; mem[2466]='h03a6; mem[2467]='h03c6; mem[2468]='h03e6; mem[2469]='h0405; mem[2470]='h0445; mem[2471]='h0485; // address 0x1340
    mem[2472]='h04c5; mem[2473]='h0505; mem[2474]='h0545; mem[2475]='h0585; mem[2476]='h05c5; mem[2477]='h0605; mem[2478]='h0645; mem[2479]='h0685; // address 0x1350
    mem[2480]='h06c5; mem[2481]='h0705; mem[2482]='h0745; mem[2483]='h0804; mem[2484]='h0904; mem[2485]='h0a04; mem[2486]='h0b04; mem[2487]='h1001; // address 0x1360
    mem[2488]='h1101; mem[2489]='h1201; mem[2490]='h1301; mem[2491]='h1401; mem[2492]='h1501; mem[2493]='h1601; mem[2494]='h1701; mem[2495]='h1801; // address 0x1370
    mem[2496]='h1901; mem[2497]='h1a01; mem[2498]='h1b01; mem[2499]='h1c01; mem[2500]='h1d09; mem[2501]='h1e09; mem[2502]='h1f09; mem[2503]='h2002; // address 0x1380
    mem[2504]='h2402; mem[2505]='h2802; mem[2506]='h2c03; mem[2507]='h3003; mem[2508]='h3403; mem[2509]='h3808; mem[2510]='h3c08; mem[2511]='h4000; // address 0x1390
    mem[2512]='h5000; mem[2513]='h6000; mem[2514]='h7000; mem[2515]='h8000; mem[2516]='h9000; mem[2517]='ha000; mem[2518]='hb000; mem[2519]='hc000; // address 0x13a0
    mem[2520]='hd000; mem[2521]='he000; mem[2522]='hf000; mem[2523]='h4c53; mem[2524]='h5420; mem[2525]='h4c57; mem[2526]='h5020; mem[2527]='h4449; // address 0x13b0
    mem[2528]='h5653; mem[2529]='h4d50; mem[2530]='h5953; mem[2531]='h4c49; mem[2532]='h2020; mem[2533]='h4149; mem[2534]='h2020; mem[2535]='h414e; // address 0x13c0
    mem[2536]='h4449; mem[2537]='h4f52; mem[2538]='h4920; mem[2539]='h4349; mem[2540]='h2020; mem[2541]='h5354; mem[2542]='h5750; mem[2543]='h5354; // address 0x13d0
    mem[2544]='h5354; mem[2545]='h4c57; mem[2546]='h5049; mem[2547]='h4c49; mem[2548]='h4d49; mem[2549]='h4944; mem[2550]='h4c45; mem[2551]='h5253; // address 0x13e0
    mem[2552]='h4554; mem[2553]='h5254; mem[2554]='h5750; mem[2555]='h434b; mem[2556]='h4f4e; mem[2557]='h434b; mem[2558]='h4f46; mem[2559]='h4c52; // address 0x13f0
    mem[2560]='h4558; mem[2561]='h424c; mem[2562]='h5750; mem[2563]='h4220; mem[2564]='h2020; mem[2565]='h5820; mem[2566]='h2020; mem[2567]='h434c; // address 0x1400
    mem[2568]='h5220; mem[2569]='h4e45; mem[2570]='h4720; mem[2571]='h494e; mem[2572]='h5620; mem[2573]='h494e; mem[2574]='h4320; mem[2575]='h494e; // address 0x1410
    mem[2576]='h4354; mem[2577]='h4445; mem[2578]='h4320; mem[2579]='h4445; mem[2580]='h4354; mem[2581]='h424c; mem[2582]='h2020; mem[2583]='h5357; // address 0x1420
    mem[2584]='h5042; mem[2585]='h5345; mem[2586]='h544f; mem[2587]='h4142; mem[2588]='h5320; mem[2589]='h5352; mem[2590]='h4120; mem[2591]='h5352; // address 0x1430
    mem[2592]='h4c20; mem[2593]='h534c; mem[2594]='h4120; mem[2595]='h5352; mem[2596]='h4320; mem[2597]='h4a4d; mem[2598]='h5020; mem[2599]='h4a4c; // address 0x1440
    mem[2600]='h5420; mem[2601]='h4a4c; mem[2602]='h4520; mem[2603]='h4a45; mem[2604]='h5120; mem[2605]='h4a48; mem[2606]='h4520; mem[2607]='h4a47; // address 0x1450
    mem[2608]='h5420; mem[2609]='h4a4e; mem[2610]='h4520; mem[2611]='h4a4e; mem[2612]='h4320; mem[2613]='h4a4f; mem[2614]='h4320; mem[2615]='h4a4e; // address 0x1460
    mem[2616]='h4f20; mem[2617]='h4a4c; mem[2618]='h2020; mem[2619]='h4a48; mem[2620]='h2020; mem[2621]='h4a4f; mem[2622]='h5020; mem[2623]='h5342; // address 0x1470
    mem[2624]='h4f20; mem[2625]='h5342; mem[2626]='h5a20; mem[2627]='h5442; mem[2628]='h2020; mem[2629]='h434f; mem[2630]='h4320; mem[2631]='h435a; // address 0x1480
    mem[2632]='h4320; mem[2633]='h584f; mem[2634]='h5220; mem[2635]='h584f; mem[2636]='h5020; mem[2637]='h4c44; mem[2638]='h4352; mem[2639]='h5354; // address 0x1490
    mem[2640]='h4352; mem[2641]='h4d50; mem[2642]='h5920; mem[2643]='h4449; mem[2644]='h5620; mem[2645]='h535a; mem[2646]='h4320; mem[2647]='h535a; // address 0x14a0
    mem[2648]='h4342; mem[2649]='h5320; mem[2650]='h2020; mem[2651]='h5342; mem[2652]='h2020; mem[2653]='h4320; mem[2654]='h2020; mem[2655]='h4342; // address 0x14b0
    mem[2656]='h2020; mem[2657]='h4120; mem[2658]='h2020; mem[2659]='h4142; mem[2660]='h2020; mem[2661]='h4d4f; mem[2662]='h5620; mem[2663]='h4d4f; // address 0x14c0
    mem[2664]='h5642; mem[2665]='h534f; mem[2666]='h4320; mem[2667]='h534f; mem[2668]='h4342; mem[2669]='h4e4f; mem[2670]='h5020; mem[2671]='h4441; // address 0x14d0
    mem[2672]='h5441; mem[2673]='h5445; mem[2674]='h5854; mem[2675]='h414f; mem[2676]='h5247; mem[2677]='h454e; mem[2678]='h4420; mem[2679]='h5254; // address 0x14e0
    mem[2680]='h2020; mem[2681]='h0000; mem[2682]='h403e; mem[2683]='h002a; mem[2684]='h5200; mem[2685]='hffff; mem[2686]='hffff; mem[2687]='hffff; // address 0x14f0
    mem[2688]='hffff; mem[2689]='hffff; mem[2690]='hffff; mem[2691]='hffff; mem[2692]='hffff; mem[2693]='hffff; mem[2694]='hffff; mem[2695]='hffff; // address 0x1500
    mem[2696]='hffff; mem[2697]='hffff; mem[2698]='hffff; mem[2699]='hffff; mem[2700]='hffff; mem[2701]='hffff; mem[2702]='hffff; mem[2703]='hffff; // address 0x1510
    mem[2704]='hffff; mem[2705]='hffff; mem[2706]='hffff; mem[2707]='hffff; mem[2708]='hffff; mem[2709]='hffff; mem[2710]='hffff; mem[2711]='hffff; // address 0x1520
    mem[2712]='hffff; mem[2713]='hffff; mem[2714]='hffff; mem[2715]='hffff; mem[2716]='hffff; mem[2717]='hffff; mem[2718]='hffff; mem[2719]='hffff; // address 0x1530
    mem[2720]='hffff; mem[2721]='hffff; mem[2722]='hffff; mem[2723]='hffff; mem[2724]='hffff; mem[2725]='hffff; mem[2726]='hffff; mem[2727]='hffff; // address 0x1540
    mem[2728]='hffff; mem[2729]='hffff; mem[2730]='hffff; mem[2731]='hffff; mem[2732]='hffff; mem[2733]='hffff; mem[2734]='hffff; mem[2735]='hffff; // address 0x1550
    mem[2736]='hffff; mem[2737]='hffff; mem[2738]='hffff; mem[2739]='hffff; mem[2740]='hffff; mem[2741]='hffff; mem[2742]='hffff; mem[2743]='hffff; // address 0x1560
    mem[2744]='hffff; mem[2745]='hffff; mem[2746]='hffff; mem[2747]='hffff; mem[2748]='hffff; mem[2749]='hffff; mem[2750]='hffff; mem[2751]='hffff; // address 0x1570
    mem[2752]='hffff; mem[2753]='hffff; mem[2754]='hffff; mem[2755]='hffff; mem[2756]='hffff; mem[2757]='hffff; mem[2758]='hffff; mem[2759]='hffff; // address 0x1580
    mem[2760]='hffff; mem[2761]='hffff; mem[2762]='hffff; mem[2763]='hffff; mem[2764]='hffff; mem[2765]='hffff; mem[2766]='hffff; mem[2767]='hffff; // address 0x1590
    mem[2768]='hffff; mem[2769]='hffff; mem[2770]='hffff; mem[2771]='hffff; mem[2772]='hffff; mem[2773]='hffff; mem[2774]='hffff; mem[2775]='hffff; // address 0x15a0
    mem[2776]='hffff; mem[2777]='hffff; mem[2778]='hffff; mem[2779]='hffff; mem[2780]='hffff; mem[2781]='hffff; mem[2782]='hffff; mem[2783]='hffff; // address 0x15b0
    mem[2784]='hffff; mem[2785]='hffff; mem[2786]='hffff; mem[2787]='hffff; mem[2788]='hffff; mem[2789]='hffff; mem[2790]='hffff; mem[2791]='hffff; // address 0x15c0
    mem[2792]='hffff; mem[2793]='hffff; mem[2794]='hffff; mem[2795]='hffff; mem[2796]='hffff; mem[2797]='hffff; mem[2798]='hffff; mem[2799]='hffff; // address 0x15d0
    mem[2800]='hffff; mem[2801]='hffff; mem[2802]='hffff; mem[2803]='hffff; mem[2804]='hffff; mem[2805]='hffff; mem[2806]='hffff; mem[2807]='hffff; // address 0x15e0
    mem[2808]='hffff; mem[2809]='hffff; mem[2810]='hffff; mem[2811]='hffff; mem[2812]='hffff; mem[2813]='hffff; mem[2814]='hffff; mem[2815]='hffff; // address 0x15f0
    mem[2816]='hffff; mem[2817]='hffff; mem[2818]='hffff; mem[2819]='hffff; mem[2820]='hffff; mem[2821]='hffff; mem[2822]='hffff; mem[2823]='hffff; // address 0x1600
    mem[2824]='hffff; mem[2825]='hffff; mem[2826]='hffff; mem[2827]='hffff; mem[2828]='hffff; mem[2829]='hffff; mem[2830]='hffff; mem[2831]='hffff; // address 0x1610
    mem[2832]='hffff; mem[2833]='hffff; mem[2834]='hffff; mem[2835]='hffff; mem[2836]='hffff; mem[2837]='hffff; mem[2838]='hffff; mem[2839]='hffff; // address 0x1620
    mem[2840]='hffff; mem[2841]='hffff; mem[2842]='hffff; mem[2843]='hffff; mem[2844]='hffff; mem[2845]='hffff; mem[2846]='hffff; mem[2847]='hffff; // address 0x1630
    mem[2848]='hffff; mem[2849]='hffff; mem[2850]='hffff; mem[2851]='hffff; mem[2852]='hffff; mem[2853]='hffff; mem[2854]='hffff; mem[2855]='hffff; // address 0x1640
    mem[2856]='hffff; mem[2857]='hffff; mem[2858]='hffff; mem[2859]='hffff; mem[2860]='hffff; mem[2861]='hffff; mem[2862]='hffff; mem[2863]='hffff; // address 0x1650
    mem[2864]='hffff; mem[2865]='hffff; mem[2866]='hffff; mem[2867]='hffff; mem[2868]='hffff; mem[2869]='hffff; mem[2870]='hffff; mem[2871]='hffff; // address 0x1660
    mem[2872]='hffff; mem[2873]='hffff; mem[2874]='hffff; mem[2875]='hffff; mem[2876]='hffff; mem[2877]='hffff; mem[2878]='hffff; mem[2879]='hffff; // address 0x1670
    mem[2880]='hffff; mem[2881]='hffff; mem[2882]='hffff; mem[2883]='hffff; mem[2884]='hffff; mem[2885]='hffff; mem[2886]='hffff; mem[2887]='hffff; // address 0x1680
    mem[2888]='hffff; mem[2889]='hffff; mem[2890]='hffff; mem[2891]='hffff; mem[2892]='hffff; mem[2893]='hffff; mem[2894]='hffff; mem[2895]='hffff; // address 0x1690
    mem[2896]='hffff; mem[2897]='hffff; mem[2898]='hffff; mem[2899]='hffff; mem[2900]='hffff; mem[2901]='hffff; mem[2902]='hffff; mem[2903]='hffff; // address 0x16a0
    mem[2904]='hffff; mem[2905]='hffff; mem[2906]='hffff; mem[2907]='hffff; mem[2908]='hffff; mem[2909]='hffff; mem[2910]='hffff; mem[2911]='hffff; // address 0x16b0
    mem[2912]='hffff; mem[2913]='hffff; mem[2914]='hffff; mem[2915]='hffff; mem[2916]='hffff; mem[2917]='hffff; mem[2918]='hffff; mem[2919]='hffff; // address 0x16c0
    mem[2920]='hffff; mem[2921]='hffff; mem[2922]='hffff; mem[2923]='hffff; mem[2924]='hffff; mem[2925]='hffff; mem[2926]='hffff; mem[2927]='hffff; // address 0x16d0
    mem[2928]='hffff; mem[2929]='hffff; mem[2930]='hffff; mem[2931]='hffff; mem[2932]='hffff; mem[2933]='hffff; mem[2934]='hffff; mem[2935]='hffff; // address 0x16e0
    mem[2936]='hffff; mem[2937]='hffff; mem[2938]='hffff; mem[2939]='hffff; mem[2940]='hffff; mem[2941]='hffff; mem[2942]='hffff; mem[2943]='hffff; // address 0x16f0
    mem[2944]='hffff; mem[2945]='hffff; mem[2946]='hffff; mem[2947]='hffff; mem[2948]='hffff; mem[2949]='hffff; mem[2950]='hffff; mem[2951]='hffff; // address 0x1700
    mem[2952]='hffff; mem[2953]='hffff; mem[2954]='hffff; mem[2955]='hffff; mem[2956]='hffff; mem[2957]='hffff; mem[2958]='hffff; mem[2959]='hffff; // address 0x1710
    mem[2960]='hffff; mem[2961]='hffff; mem[2962]='hffff; mem[2963]='hffff; mem[2964]='hffff; mem[2965]='hffff; mem[2966]='hffff; mem[2967]='hffff; // address 0x1720
    mem[2968]='hffff; mem[2969]='hffff; mem[2970]='hffff; mem[2971]='hffff; mem[2972]='hffff; mem[2973]='hffff; mem[2974]='hffff; mem[2975]='hffff; // address 0x1730
    mem[2976]='hffff; mem[2977]='hffff; mem[2978]='hffff; mem[2979]='hffff; mem[2980]='hffff; mem[2981]='hffff; mem[2982]='hffff; mem[2983]='hffff; // address 0x1740
    mem[2984]='hffff; mem[2985]='hffff; mem[2986]='hffff; mem[2987]='hffff; mem[2988]='hffff; mem[2989]='hffff; mem[2990]='hffff; mem[2991]='hffff; // address 0x1750
    mem[2992]='hffff; mem[2993]='hffff; mem[2994]='hffff; mem[2995]='hffff; mem[2996]='hffff; mem[2997]='hffff; mem[2998]='hffff; mem[2999]='hffff; // address 0x1760
    mem[3000]='hffff; mem[3001]='hffff; mem[3002]='hffff; mem[3003]='hffff; mem[3004]='hffff; mem[3005]='hffff; mem[3006]='hffff; mem[3007]='hffff; // address 0x1770
    mem[3008]='hffff; mem[3009]='hffff; mem[3010]='hffff; mem[3011]='hffff; mem[3012]='hffff; mem[3013]='hffff; mem[3014]='hffff; mem[3015]='hffff; // address 0x1780
    mem[3016]='hffff; mem[3017]='hffff; mem[3018]='hffff; mem[3019]='hffff; mem[3020]='hffff; mem[3021]='hffff; mem[3022]='hffff; mem[3023]='hffff; // address 0x1790
    mem[3024]='hffff; mem[3025]='hffff; mem[3026]='hffff; mem[3027]='hffff; mem[3028]='hffff; mem[3029]='hffff; mem[3030]='hffff; mem[3031]='hffff; // address 0x17a0
    mem[3032]='hffff; mem[3033]='hffff; mem[3034]='hffff; mem[3035]='hffff; mem[3036]='hffff; mem[3037]='hffff; mem[3038]='hffff; mem[3039]='hffff; // address 0x17b0
    mem[3040]='hffff; mem[3041]='hffff; mem[3042]='hffff; mem[3043]='hffff; mem[3044]='hffff; mem[3045]='hffff; mem[3046]='hffff; mem[3047]='hffff; // address 0x17c0
    mem[3048]='hffff; mem[3049]='hffff; mem[3050]='hffff; mem[3051]='hffff; mem[3052]='hffff; mem[3053]='hffff; mem[3054]='hffff; mem[3055]='hffff; // address 0x17d0
    mem[3056]='hffff; mem[3057]='hffff; mem[3058]='hffff; mem[3059]='hffff; mem[3060]='hffff; mem[3061]='hffff; mem[3062]='hffff; mem[3063]='hffff; // address 0x17e0
    mem[3064]='hffff; mem[3065]='hffff; mem[3066]='hffff; mem[3067]='hffff; mem[3068]='hffff; mem[3069]='hffff; mem[3070]='hffff; mem[3071]='hffff; // address 0x17f0
    mem[3072]='hffff; mem[3073]='hffff; mem[3074]='hffff; mem[3075]='hffff; mem[3076]='hffff; mem[3077]='hffff; mem[3078]='hffff; mem[3079]='hffff; // address 0x1800
    mem[3080]='hffff; mem[3081]='hffff; mem[3082]='hffff; mem[3083]='hffff; mem[3084]='hffff; mem[3085]='hffff; mem[3086]='hffff; mem[3087]='hffff; // address 0x1810
    mem[3088]='hffff; mem[3089]='hffff; mem[3090]='hffff; mem[3091]='hffff; mem[3092]='hffff; mem[3093]='hffff; mem[3094]='hffff; mem[3095]='hffff; // address 0x1820
    mem[3096]='hffff; mem[3097]='hffff; mem[3098]='hffff; mem[3099]='hffff; mem[3100]='hffff; mem[3101]='hffff; mem[3102]='hffff; mem[3103]='hffff; // address 0x1830
    mem[3104]='hffff; mem[3105]='hffff; mem[3106]='hffff; mem[3107]='hffff; mem[3108]='hffff; mem[3109]='hffff; mem[3110]='hffff; mem[3111]='hffff; // address 0x1840
    mem[3112]='hffff; mem[3113]='hffff; mem[3114]='hffff; mem[3115]='hffff; mem[3116]='hffff; mem[3117]='hffff; mem[3118]='hffff; mem[3119]='hffff; // address 0x1850
    mem[3120]='hffff; mem[3121]='hffff; mem[3122]='hffff; mem[3123]='hffff; mem[3124]='hffff; mem[3125]='hffff; mem[3126]='hffff; mem[3127]='hffff; // address 0x1860
    mem[3128]='hffff; mem[3129]='hffff; mem[3130]='hffff; mem[3131]='hffff; mem[3132]='hffff; mem[3133]='hffff; mem[3134]='hffff; mem[3135]='hffff; // address 0x1870
    mem[3136]='hffff; mem[3137]='hffff; mem[3138]='hffff; mem[3139]='hffff; mem[3140]='hffff; mem[3141]='hffff; mem[3142]='hffff; mem[3143]='hffff; // address 0x1880
    mem[3144]='hffff; mem[3145]='hffff; mem[3146]='hffff; mem[3147]='hffff; mem[3148]='hffff; mem[3149]='hffff; mem[3150]='hffff; mem[3151]='hffff; // address 0x1890
    mem[3152]='hffff; mem[3153]='hffff; mem[3154]='hffff; mem[3155]='hffff; mem[3156]='hffff; mem[3157]='hffff; mem[3158]='hffff; mem[3159]='hffff; // address 0x18a0
    mem[3160]='hffff; mem[3161]='hffff; mem[3162]='hffff; mem[3163]='hffff; mem[3164]='hffff; mem[3165]='hffff; mem[3166]='hffff; mem[3167]='hffff; // address 0x18b0
    mem[3168]='hffff; mem[3169]='hffff; mem[3170]='hffff; mem[3171]='hffff; mem[3172]='hffff; mem[3173]='hffff; mem[3174]='hffff; mem[3175]='hffff; // address 0x18c0
    mem[3176]='hffff; mem[3177]='hffff; mem[3178]='hffff; mem[3179]='hffff; mem[3180]='hffff; mem[3181]='hffff; mem[3182]='hffff; mem[3183]='hffff; // address 0x18d0
    mem[3184]='hffff; mem[3185]='hffff; mem[3186]='hffff; mem[3187]='hffff; mem[3188]='hffff; mem[3189]='hffff; mem[3190]='hffff; mem[3191]='hffff; // address 0x18e0
    mem[3192]='hffff; mem[3193]='hffff; mem[3194]='hffff; mem[3195]='hffff; mem[3196]='hffff; mem[3197]='hffff; mem[3198]='hffff; mem[3199]='hffff; // address 0x18f0
    mem[3200]='hffff; mem[3201]='hffff; mem[3202]='hffff; mem[3203]='hffff; mem[3204]='hffff; mem[3205]='hffff; mem[3206]='hffff; mem[3207]='hffff; // address 0x1900
    mem[3208]='hffff; mem[3209]='hffff; mem[3210]='hffff; mem[3211]='hffff; mem[3212]='hffff; mem[3213]='hffff; mem[3214]='hffff; mem[3215]='hffff; // address 0x1910
    mem[3216]='hffff; mem[3217]='hffff; mem[3218]='hffff; mem[3219]='hffff; mem[3220]='hffff; mem[3221]='hffff; mem[3222]='hffff; mem[3223]='hffff; // address 0x1920
    mem[3224]='hffff; mem[3225]='hffff; mem[3226]='hffff; mem[3227]='hffff; mem[3228]='hffff; mem[3229]='hffff; mem[3230]='hffff; mem[3231]='hffff; // address 0x1930
    mem[3232]='hffff; mem[3233]='hffff; mem[3234]='hffff; mem[3235]='hffff; mem[3236]='hffff; mem[3237]='hffff; mem[3238]='hffff; mem[3239]='hffff; // address 0x1940
    mem[3240]='hffff; mem[3241]='hffff; mem[3242]='hffff; mem[3243]='hffff; mem[3244]='hffff; mem[3245]='hffff; mem[3246]='hffff; mem[3247]='hffff; // address 0x1950
    mem[3248]='hffff; mem[3249]='hffff; mem[3250]='hffff; mem[3251]='hffff; mem[3252]='hffff; mem[3253]='hffff; mem[3254]='hffff; mem[3255]='hffff; // address 0x1960
    mem[3256]='hffff; mem[3257]='hffff; mem[3258]='hffff; mem[3259]='hffff; mem[3260]='hffff; mem[3261]='hffff; mem[3262]='hffff; mem[3263]='hffff; // address 0x1970
    mem[3264]='hffff; mem[3265]='hffff; mem[3266]='hffff; mem[3267]='hffff; mem[3268]='hffff; mem[3269]='hffff; mem[3270]='hffff; mem[3271]='hffff; // address 0x1980
    mem[3272]='hffff; mem[3273]='hffff; mem[3274]='hffff; mem[3275]='hffff; mem[3276]='hffff; mem[3277]='hffff; mem[3278]='hffff; mem[3279]='hffff; // address 0x1990
    mem[3280]='hffff; mem[3281]='hffff; mem[3282]='hffff; mem[3283]='hffff; mem[3284]='hffff; mem[3285]='hffff; mem[3286]='hffff; mem[3287]='hffff; // address 0x19a0
    mem[3288]='hffff; mem[3289]='hffff; mem[3290]='hffff; mem[3291]='hffff; mem[3292]='hffff; mem[3293]='hffff; mem[3294]='hffff; mem[3295]='hffff; // address 0x19b0
    mem[3296]='hffff; mem[3297]='hffff; mem[3298]='hffff; mem[3299]='hffff; mem[3300]='hffff; mem[3301]='hffff; mem[3302]='hffff; mem[3303]='hffff; // address 0x19c0
    mem[3304]='hffff; mem[3305]='hffff; mem[3306]='hffff; mem[3307]='hffff; mem[3308]='hffff; mem[3309]='hffff; mem[3310]='hffff; mem[3311]='hffff; // address 0x19d0
    mem[3312]='hffff; mem[3313]='hffff; mem[3314]='hffff; mem[3315]='hffff; mem[3316]='hffff; mem[3317]='hffff; mem[3318]='hffff; mem[3319]='hffff; // address 0x19e0
    mem[3320]='hffff; mem[3321]='hffff; mem[3322]='hffff; mem[3323]='hffff; mem[3324]='hffff; mem[3325]='hffff; mem[3326]='hffff; mem[3327]='hffff; // address 0x19f0
    mem[3328]='hffff; mem[3329]='hffff; mem[3330]='hffff; mem[3331]='hffff; mem[3332]='hffff; mem[3333]='hffff; mem[3334]='hffff; mem[3335]='hffff; // address 0x1a00
    mem[3336]='hffff; mem[3337]='hffff; mem[3338]='hffff; mem[3339]='hffff; mem[3340]='hffff; mem[3341]='hffff; mem[3342]='hffff; mem[3343]='hffff; // address 0x1a10
    mem[3344]='hffff; mem[3345]='hffff; mem[3346]='hffff; mem[3347]='hffff; mem[3348]='hffff; mem[3349]='hffff; mem[3350]='hffff; mem[3351]='hffff; // address 0x1a20
    mem[3352]='hffff; mem[3353]='hffff; mem[3354]='hffff; mem[3355]='hffff; mem[3356]='hffff; mem[3357]='hffff; mem[3358]='hffff; mem[3359]='hffff; // address 0x1a30
    mem[3360]='hffff; mem[3361]='hffff; mem[3362]='hffff; mem[3363]='hffff; mem[3364]='hffff; mem[3365]='hffff; mem[3366]='hffff; mem[3367]='hffff; // address 0x1a40
    mem[3368]='hffff; mem[3369]='hffff; mem[3370]='hffff; mem[3371]='hffff; mem[3372]='hffff; mem[3373]='hffff; mem[3374]='hffff; mem[3375]='hffff; // address 0x1a50
    mem[3376]='hffff; mem[3377]='hffff; mem[3378]='hffff; mem[3379]='hffff; mem[3380]='hffff; mem[3381]='hffff; mem[3382]='hffff; mem[3383]='hffff; // address 0x1a60
    mem[3384]='hffff; mem[3385]='hffff; mem[3386]='hffff; mem[3387]='hffff; mem[3388]='hffff; mem[3389]='hffff; mem[3390]='hffff; mem[3391]='hffff; // address 0x1a70
    mem[3392]='hffff; mem[3393]='hffff; mem[3394]='hffff; mem[3395]='hffff; mem[3396]='hffff; mem[3397]='hffff; mem[3398]='hffff; mem[3399]='hffff; // address 0x1a80
    mem[3400]='hffff; mem[3401]='hffff; mem[3402]='hffff; mem[3403]='hffff; mem[3404]='hffff; mem[3405]='hffff; mem[3406]='hffff; mem[3407]='hffff; // address 0x1a90
    mem[3408]='hffff; mem[3409]='hffff; mem[3410]='hffff; mem[3411]='hffff; mem[3412]='hffff; mem[3413]='hffff; mem[3414]='hffff; mem[3415]='hffff; // address 0x1aa0
    mem[3416]='hffff; mem[3417]='hffff; mem[3418]='hffff; mem[3419]='hffff; mem[3420]='hffff; mem[3421]='hffff; mem[3422]='hffff; mem[3423]='hffff; // address 0x1ab0
    mem[3424]='hffff; mem[3425]='hffff; mem[3426]='hffff; mem[3427]='hffff; mem[3428]='hffff; mem[3429]='hffff; mem[3430]='hffff; mem[3431]='hffff; // address 0x1ac0
    mem[3432]='hffff; mem[3433]='hffff; mem[3434]='hffff; mem[3435]='hffff; mem[3436]='hffff; mem[3437]='hffff; mem[3438]='hffff; mem[3439]='hffff; // address 0x1ad0
    mem[3440]='hffff; mem[3441]='hffff; mem[3442]='hffff; mem[3443]='hffff; mem[3444]='hffff; mem[3445]='hffff; mem[3446]='hffff; mem[3447]='hffff; // address 0x1ae0
    mem[3448]='hffff; mem[3449]='hffff; mem[3450]='hffff; mem[3451]='hffff; mem[3452]='hffff; mem[3453]='hffff; mem[3454]='hffff; mem[3455]='hffff; // address 0x1af0
    mem[3456]='hffff; mem[3457]='hffff; mem[3458]='hffff; mem[3459]='hffff; mem[3460]='hffff; mem[3461]='hffff; mem[3462]='hffff; mem[3463]='hffff; // address 0x1b00
    mem[3464]='hffff; mem[3465]='hffff; mem[3466]='hffff; mem[3467]='hffff; mem[3468]='hffff; mem[3469]='hffff; mem[3470]='hffff; mem[3471]='hffff; // address 0x1b10
    mem[3472]='hffff; mem[3473]='hffff; mem[3474]='hffff; mem[3475]='hffff; mem[3476]='hffff; mem[3477]='hffff; mem[3478]='hffff; mem[3479]='hffff; // address 0x1b20
    mem[3480]='hffff; mem[3481]='hffff; mem[3482]='hffff; mem[3483]='hffff; mem[3484]='hffff; mem[3485]='hffff; mem[3486]='hffff; mem[3487]='hffff; // address 0x1b30
    mem[3488]='hffff; mem[3489]='hffff; mem[3490]='hffff; mem[3491]='hffff; mem[3492]='hffff; mem[3493]='hffff; mem[3494]='hffff; mem[3495]='hffff; // address 0x1b40
    mem[3496]='hffff; mem[3497]='hffff; mem[3498]='hffff; mem[3499]='hffff; mem[3500]='hffff; mem[3501]='hffff; mem[3502]='hffff; mem[3503]='hffff; // address 0x1b50
    mem[3504]='hffff; mem[3505]='hffff; mem[3506]='hffff; mem[3507]='hffff; mem[3508]='hffff; mem[3509]='hffff; mem[3510]='hffff; mem[3511]='hffff; // address 0x1b60
    mem[3512]='hffff; mem[3513]='hffff; mem[3514]='hffff; mem[3515]='hffff; mem[3516]='hffff; mem[3517]='hffff; mem[3518]='hffff; mem[3519]='hffff; // address 0x1b70
    mem[3520]='hffff; mem[3521]='hffff; mem[3522]='hffff; mem[3523]='hffff; mem[3524]='hffff; mem[3525]='hffff; mem[3526]='hffff; mem[3527]='hffff; // address 0x1b80
    mem[3528]='hffff; mem[3529]='hffff; mem[3530]='hffff; mem[3531]='hffff; mem[3532]='hffff; mem[3533]='hffff; mem[3534]='hffff; mem[3535]='hffff; // address 0x1b90
    mem[3536]='hffff; mem[3537]='hffff; mem[3538]='hffff; mem[3539]='hffff; mem[3540]='hffff; mem[3541]='hffff; mem[3542]='hffff; mem[3543]='hffff; // address 0x1ba0
    mem[3544]='hffff; mem[3545]='hffff; mem[3546]='hffff; mem[3547]='hffff; mem[3548]='hffff; mem[3549]='hffff; mem[3550]='hffff; mem[3551]='hffff; // address 0x1bb0
    mem[3552]='hffff; mem[3553]='hffff; mem[3554]='hffff; mem[3555]='hffff; mem[3556]='hffff; mem[3557]='hffff; mem[3558]='hffff; mem[3559]='hffff; // address 0x1bc0
    mem[3560]='hffff; mem[3561]='hffff; mem[3562]='hffff; mem[3563]='hffff; mem[3564]='hffff; mem[3565]='hffff; mem[3566]='hffff; mem[3567]='hffff; // address 0x1bd0
    mem[3568]='hffff; mem[3569]='hffff; mem[3570]='hffff; mem[3571]='hffff; mem[3572]='hffff; mem[3573]='hffff; mem[3574]='hffff; mem[3575]='hffff; // address 0x1be0
    mem[3576]='hffff; mem[3577]='hffff; mem[3578]='hffff; mem[3579]='hffff; mem[3580]='hffff; mem[3581]='hffff; mem[3582]='hffff; mem[3583]='hffff; // address 0x1bf0
    mem[3584]='hffff; mem[3585]='hffff; mem[3586]='hffff; mem[3587]='hffff; mem[3588]='hffff; mem[3589]='hffff; mem[3590]='hffff; mem[3591]='hffff; // address 0x1c00
    mem[3592]='hffff; mem[3593]='hffff; mem[3594]='hffff; mem[3595]='hffff; mem[3596]='hffff; mem[3597]='hffff; mem[3598]='hffff; mem[3599]='hffff; // address 0x1c10
    mem[3600]='hffff; mem[3601]='hffff; mem[3602]='hffff; mem[3603]='hffff; mem[3604]='hffff; mem[3605]='hffff; mem[3606]='hffff; mem[3607]='hffff; // address 0x1c20
    mem[3608]='hffff; mem[3609]='hffff; mem[3610]='hffff; mem[3611]='hffff; mem[3612]='hffff; mem[3613]='hffff; mem[3614]='hffff; mem[3615]='hffff; // address 0x1c30
    mem[3616]='hffff; mem[3617]='hffff; mem[3618]='hffff; mem[3619]='hffff; mem[3620]='hffff; mem[3621]='hffff; mem[3622]='hffff; mem[3623]='hffff; // address 0x1c40
    mem[3624]='hffff; mem[3625]='hffff; mem[3626]='hffff; mem[3627]='hffff; mem[3628]='hffff; mem[3629]='hffff; mem[3630]='hffff; mem[3631]='hffff; // address 0x1c50
    mem[3632]='hffff; mem[3633]='hffff; mem[3634]='hffff; mem[3635]='hffff; mem[3636]='hffff; mem[3637]='hffff; mem[3638]='hffff; mem[3639]='hffff; // address 0x1c60
    mem[3640]='hffff; mem[3641]='hffff; mem[3642]='hffff; mem[3643]='hffff; mem[3644]='hffff; mem[3645]='hffff; mem[3646]='hffff; mem[3647]='hffff; // address 0x1c70
    mem[3648]='hffff; mem[3649]='hffff; mem[3650]='hffff; mem[3651]='hffff; mem[3652]='hffff; mem[3653]='hffff; mem[3654]='hffff; mem[3655]='hffff; // address 0x1c80
    mem[3656]='hffff; mem[3657]='hffff; mem[3658]='hffff; mem[3659]='hffff; mem[3660]='hffff; mem[3661]='hffff; mem[3662]='hffff; mem[3663]='hffff; // address 0x1c90
    mem[3664]='hffff; mem[3665]='hffff; mem[3666]='hffff; mem[3667]='hffff; mem[3668]='hffff; mem[3669]='hffff; mem[3670]='hffff; mem[3671]='hffff; // address 0x1ca0
    mem[3672]='hffff; mem[3673]='hffff; mem[3674]='hffff; mem[3675]='hffff; mem[3676]='hffff; mem[3677]='hffff; mem[3678]='hffff; mem[3679]='hffff; // address 0x1cb0
    mem[3680]='hffff; mem[3681]='hffff; mem[3682]='hffff; mem[3683]='hffff; mem[3684]='hffff; mem[3685]='hffff; mem[3686]='hffff; mem[3687]='hffff; // address 0x1cc0
    mem[3688]='hffff; mem[3689]='hffff; mem[3690]='hffff; mem[3691]='hffff; mem[3692]='hffff; mem[3693]='hffff; mem[3694]='hffff; mem[3695]='hffff; // address 0x1cd0
    mem[3696]='hffff; mem[3697]='hffff; mem[3698]='hffff; mem[3699]='hffff; mem[3700]='hffff; mem[3701]='hffff; mem[3702]='hffff; mem[3703]='hffff; // address 0x1ce0
    mem[3704]='hffff; mem[3705]='hffff; mem[3706]='hffff; mem[3707]='hffff; mem[3708]='hffff; mem[3709]='hffff; mem[3710]='hffff; mem[3711]='hffff; // address 0x1cf0
    mem[3712]='hffff; mem[3713]='hffff; mem[3714]='hffff; mem[3715]='hffff; mem[3716]='hffff; mem[3717]='hffff; mem[3718]='hffff; mem[3719]='hffff; // address 0x1d00
    mem[3720]='hffff; mem[3721]='hffff; mem[3722]='hffff; mem[3723]='hffff; mem[3724]='hffff; mem[3725]='hffff; mem[3726]='hffff; mem[3727]='hffff; // address 0x1d10
    mem[3728]='hffff; mem[3729]='hffff; mem[3730]='hffff; mem[3731]='hffff; mem[3732]='hffff; mem[3733]='hffff; mem[3734]='hffff; mem[3735]='hffff; // address 0x1d20
    mem[3736]='hffff; mem[3737]='hffff; mem[3738]='hffff; mem[3739]='hffff; mem[3740]='hffff; mem[3741]='hffff; mem[3742]='hffff; mem[3743]='hffff; // address 0x1d30
    mem[3744]='hffff; mem[3745]='hffff; mem[3746]='hffff; mem[3747]='hffff; mem[3748]='hffff; mem[3749]='hffff; mem[3750]='hffff; mem[3751]='hffff; // address 0x1d40
    mem[3752]='hffff; mem[3753]='hffff; mem[3754]='hffff; mem[3755]='hffff; mem[3756]='hffff; mem[3757]='hffff; mem[3758]='hffff; mem[3759]='hffff; // address 0x1d50
    mem[3760]='hffff; mem[3761]='hffff; mem[3762]='hffff; mem[3763]='hffff; mem[3764]='hffff; mem[3765]='hffff; mem[3766]='hffff; mem[3767]='hffff; // address 0x1d60
    mem[3768]='hffff; mem[3769]='hffff; mem[3770]='hffff; mem[3771]='hffff; mem[3772]='hffff; mem[3773]='hffff; mem[3774]='hffff; mem[3775]='hffff; // address 0x1d70
    mem[3776]='hffff; mem[3777]='hffff; mem[3778]='hffff; mem[3779]='hffff; mem[3780]='hffff; mem[3781]='hffff; mem[3782]='hffff; mem[3783]='hffff; // address 0x1d80
    mem[3784]='hffff; mem[3785]='hffff; mem[3786]='hffff; mem[3787]='hffff; mem[3788]='hffff; mem[3789]='hffff; mem[3790]='hffff; mem[3791]='hffff; // address 0x1d90
    mem[3792]='hffff; mem[3793]='hffff; mem[3794]='hffff; mem[3795]='hffff; mem[3796]='hffff; mem[3797]='hffff; mem[3798]='hffff; mem[3799]='hffff; // address 0x1da0
    mem[3800]='hffff; mem[3801]='hffff; mem[3802]='hffff; mem[3803]='hffff; mem[3804]='hffff; mem[3805]='hffff; mem[3806]='hffff; mem[3807]='hffff; // address 0x1db0
    mem[3808]='hffff; mem[3809]='hffff; mem[3810]='hffff; mem[3811]='hffff; mem[3812]='hffff; mem[3813]='hffff; mem[3814]='hffff; mem[3815]='hffff; // address 0x1dc0
    mem[3816]='hffff; mem[3817]='hffff; mem[3818]='hffff; mem[3819]='hffff; mem[3820]='hffff; mem[3821]='hffff; mem[3822]='hffff; mem[3823]='hffff; // address 0x1dd0
    mem[3824]='hffff; mem[3825]='hffff; mem[3826]='hffff; mem[3827]='hffff; mem[3828]='hffff; mem[3829]='hffff; mem[3830]='hffff; mem[3831]='hffff; // address 0x1de0
    mem[3832]='hffff; mem[3833]='hffff; mem[3834]='hffff; mem[3835]='hffff; mem[3836]='hffff; mem[3837]='hffff; mem[3838]='hffff; mem[3839]='hffff; // address 0x1df0
    mem[3840]='hffff; mem[3841]='hffff; mem[3842]='hffff; mem[3843]='hffff; mem[3844]='hffff; mem[3845]='hffff; mem[3846]='hffff; mem[3847]='hffff; // address 0x1e00
    mem[3848]='hffff; mem[3849]='hffff; mem[3850]='hffff; mem[3851]='hffff; mem[3852]='hffff; mem[3853]='hffff; mem[3854]='hffff; mem[3855]='hffff; // address 0x1e10
    mem[3856]='hffff; mem[3857]='hffff; mem[3858]='hffff; mem[3859]='hffff; mem[3860]='hffff; mem[3861]='hffff; mem[3862]='hffff; mem[3863]='hffff; // address 0x1e20
    mem[3864]='hffff; mem[3865]='hffff; mem[3866]='hffff; mem[3867]='hffff; mem[3868]='hffff; mem[3869]='hffff; mem[3870]='hffff; mem[3871]='hffff; // address 0x1e30
    mem[3872]='hffff; mem[3873]='hffff; mem[3874]='hffff; mem[3875]='hffff; mem[3876]='hffff; mem[3877]='hffff; mem[3878]='hffff; mem[3879]='hffff; // address 0x1e40
    mem[3880]='hffff; mem[3881]='hffff; mem[3882]='hffff; mem[3883]='hffff; mem[3884]='hffff; mem[3885]='hffff; mem[3886]='hffff; mem[3887]='hffff; // address 0x1e50
    mem[3888]='hffff; mem[3889]='hffff; mem[3890]='hffff; mem[3891]='hffff; mem[3892]='hffff; mem[3893]='hffff; mem[3894]='hffff; mem[3895]='hffff; // address 0x1e60
    mem[3896]='hffff; mem[3897]='hffff; mem[3898]='hffff; mem[3899]='hffff; mem[3900]='hffff; mem[3901]='hffff; mem[3902]='hffff; mem[3903]='hffff; // address 0x1e70
    mem[3904]='hffff; mem[3905]='hffff; mem[3906]='hffff; mem[3907]='hffff; mem[3908]='hffff; mem[3909]='hffff; mem[3910]='hffff; mem[3911]='hffff; // address 0x1e80
    mem[3912]='hffff; mem[3913]='hffff; mem[3914]='hffff; mem[3915]='hffff; mem[3916]='hffff; mem[3917]='hffff; mem[3918]='hffff; mem[3919]='hffff; // address 0x1e90
    mem[3920]='hffff; mem[3921]='hffff; mem[3922]='hffff; mem[3923]='hffff; mem[3924]='hffff; mem[3925]='hffff; mem[3926]='hffff; mem[3927]='hffff; // address 0x1ea0
    mem[3928]='hffff; mem[3929]='hffff; mem[3930]='hffff; mem[3931]='hffff; mem[3932]='hffff; mem[3933]='hffff; mem[3934]='hffff; mem[3935]='hffff; // address 0x1eb0
    mem[3936]='hffff; mem[3937]='hffff; mem[3938]='hffff; mem[3939]='hffff; mem[3940]='hffff; mem[3941]='hffff; mem[3942]='hffff; mem[3943]='hffff; // address 0x1ec0
    mem[3944]='hffff; mem[3945]='hffff; mem[3946]='hffff; mem[3947]='hffff; mem[3948]='hffff; mem[3949]='hffff; mem[3950]='hffff; mem[3951]='hffff; // address 0x1ed0
    mem[3952]='hffff; mem[3953]='hffff; mem[3954]='hffff; mem[3955]='hffff; mem[3956]='hffff; mem[3957]='hffff; mem[3958]='hffff; mem[3959]='hffff; // address 0x1ee0
    mem[3960]='hffff; mem[3961]='hffff; mem[3962]='hffff; mem[3963]='hffff; mem[3964]='hffff; mem[3965]='hffff; mem[3966]='hffff; mem[3967]='hffff; // address 0x1ef0
    mem[3968]='hffff; mem[3969]='hffff; mem[3970]='hffff; mem[3971]='hffff; mem[3972]='hffff; mem[3973]='hffff; mem[3974]='hffff; mem[3975]='hffff; // address 0x1f00
    mem[3976]='hffff; mem[3977]='hffff; mem[3978]='hffff; mem[3979]='hffff; mem[3980]='hffff; mem[3981]='hffff; mem[3982]='hffff; mem[3983]='hffff; // address 0x1f10
    mem[3984]='hffff; mem[3985]='hffff; mem[3986]='hffff; mem[3987]='hffff; mem[3988]='hffff; mem[3989]='hffff; mem[3990]='hffff; mem[3991]='hffff; // address 0x1f20
    mem[3992]='hffff; mem[3993]='hffff; mem[3994]='hffff; mem[3995]='hffff; mem[3996]='hffff; mem[3997]='hffff; mem[3998]='hffff; mem[3999]='hffff; // address 0x1f30
    mem[4000]='hffff; mem[4001]='hffff; mem[4002]='hffff; mem[4003]='hffff; mem[4004]='hffff; mem[4005]='hffff; mem[4006]='hffff; mem[4007]='hffff; // address 0x1f40
    mem[4008]='hffff; mem[4009]='hffff; mem[4010]='hffff; mem[4011]='hffff; mem[4012]='hffff; mem[4013]='hffff; mem[4014]='hffff; mem[4015]='hffff; // address 0x1f50
    mem[4016]='hffff; mem[4017]='hffff; mem[4018]='hffff; mem[4019]='hffff; mem[4020]='hffff; mem[4021]='hffff; mem[4022]='hffff; mem[4023]='hffff; // address 0x1f60
    mem[4024]='hffff; mem[4025]='hffff; mem[4026]='hffff; mem[4027]='hffff; mem[4028]='hffff; mem[4029]='hffff; mem[4030]='hffff; mem[4031]='hffff; // address 0x1f70
    mem[4032]='hffff; mem[4033]='hffff; mem[4034]='hffff; mem[4035]='hffff; mem[4036]='hffff; mem[4037]='hffff; mem[4038]='hffff; mem[4039]='hffff; // address 0x1f80
    mem[4040]='hffff; mem[4041]='hffff; mem[4042]='hffff; mem[4043]='hffff; mem[4044]='hffff; mem[4045]='hffff; mem[4046]='hffff; mem[4047]='hffff; // address 0x1f90
    mem[4048]='hffff; mem[4049]='hffff; mem[4050]='hffff; mem[4051]='hffff; mem[4052]='hffff; mem[4053]='hffff; mem[4054]='hffff; mem[4055]='hffff; // address 0x1fa0
    mem[4056]='hffff; mem[4057]='hffff; mem[4058]='hffff; mem[4059]='hffff; mem[4060]='hffff; mem[4061]='hffff; mem[4062]='hffff; mem[4063]='hffff; // address 0x1fb0
    mem[4064]='hffff; mem[4065]='hffff; mem[4066]='hffff; mem[4067]='hffff; mem[4068]='hffff; mem[4069]='hffff; mem[4070]='hffff; mem[4071]='hffff; // address 0x1fc0
    mem[4072]='hffff; mem[4073]='hffff; mem[4074]='hffff; mem[4075]='hffff; mem[4076]='hffff; mem[4077]='hffff; mem[4078]='hffff; mem[4079]='hffff; // address 0x1fd0
    mem[4080]='hffff; mem[4081]='hffff; mem[4082]='hffff; mem[4083]='hffff; mem[4084]='hffff; mem[4085]='hffff; mem[4086]='hffff; mem[4087]='hffff; // address 0x1fe0
    mem[4088]='hffff; mem[4089]='hffff; mem[4090]='hffff; mem[4091]='hffff; mem[4092]='hffff; mem[4093]='hffff; mem[4094]='hffff; mem[4095]='hffff; // address 0x1ff0

    // // EP patch the ROM with test software
    // test division
    // note this breaks regular execution
/*    
    mem[4000] = 'h0202;
    mem[4001] = 'h0000; // LI R2,0
    mem[4002] = 'h0203;
    mem[4003] = 'h0064; // LI R3,100
    mem[4004] = 'h0204;
    mem[4005] = 'h0007; // LI R4,7
    mem[4006] = 'h3C84; // DIV R4,R2 = result Q=14, R=2
    mem[4007] = 'h3902; // MPY R2,R4: R4=0 (high word) R5=98
    mem[4008] = 'h0202; // LI R2,FFFF
    mem[4009] = 'hffff;
    mem[4010] = 'h0204; // LI R2,FFFF
    mem[4011] = 'hffff;
    mem[4012] = 'h3902; // MPY R2,R4: 

    mem[185] = 'h0460;  // B 8000 (decimal, hex 1f40)
    mem[186] = 'h1f40;
*/
//


    // mem[4000]='h0202; // at 8000 (1f40 hex)
    // mem[4001]='h0A05;
    // mem[4002]='h0204;
    // mem[4003]='h1234;
    // mem[4004]='h2e84;
    // mem[4005]='h0204;
    // mem[4006]='habba;

    // mem[4007]='h0202; // LI R2,>0a55 
    // mem[4008]='h0a54; // opcode for (SLA R4,5)
    // mem[4009]='h0482; // X R2

    // mem[4010]='h2e84; // XOP R4,10

    // mem[4011]='h0460; // B 0x176
    // mem[4012]='h0176;
    // // trampoline
    // mem[185]='h0460;  // B 8000 (decimal, hex 1f40)
    // mem[186]='h1f40;



  end
  
endmodule